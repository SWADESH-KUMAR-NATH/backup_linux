* SPICE3 file created from 6T-cell.ext - technology: scmos
.subckt SRAM_6T_swad q2 q1 blb bl wl example_param=1.0
M1000 q2 q1 gnd gnd scmosn w=1.2u l=0.4u
+  ad=0p pd=0u as=0p ps=0u
M1001 q1 wl bl gnd scmosn w=0.6u l=0.8u
+  ad=0p pd=0u as=0p ps=0u
M1002 q2 q1 vdd vdd scmosp w=0.6u l=1.2u
+  ad=0p pd=0u as=0p ps=0u
M1003 blb wl q2 gnd scmosn w=0.6u l=0.8u
+  ad=0p pd=0u as=0p ps=0u
M1004 vdd q2 q1 vdd scmosp w=0.6u l=1.2u
+  ad=0p pd=0u as=0p ps=0u
M1005 gnd q2 q1 gnd scmosn w=1.2u l=0.4u
+  ad=0p pd=0u as=0p ps=0u
C0 vdd q2 0.42fF
C1 q1 q2 0.42fF
C2 blb vdd 0.25fF
C3 q2 wl 0.25fF
C4 bl vdd 0.25fF
C5 blb wl 0.11fF
C6 bl q1 0.03fF
C7 q1 vdd 0.62fF
C8 bl wl 0.11fF
C9 vdd wl 0.09fF
C10 blb q2 0.03fF
C11 q1 wl 0.14fF
C12 blb gnd 0.19fF
C13 bl gnd 0.19fF
C14 wl gnd 0.79fF
C15 q1 gnd 0.29fF
C16 q2 gnd 0.45fF
C17 vdd gnd 2.86fF
.ends SRAM_6T_swad

