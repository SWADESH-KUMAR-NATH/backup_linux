magic
tech scmos
timestamp 1636204741
<< nwell >>
rect -56 22 -22 48
<< ntransistor >>
rect -44 1 -42 7
rect -36 1 -34 7
<< ptransistor >>
rect -44 28 -42 37
rect -36 28 -34 37
<< ndiffusion >>
rect -50 6 -44 7
rect -50 2 -49 6
rect -45 2 -44 6
rect -50 1 -44 2
rect -42 6 -36 7
rect -42 2 -41 6
rect -37 2 -36 6
rect -42 1 -36 2
rect -34 6 -28 7
rect -34 2 -33 6
rect -29 2 -28 6
rect -34 1 -28 2
<< pdiffusion >>
rect -50 36 -44 37
rect -50 29 -49 36
rect -45 29 -44 36
rect -50 28 -44 29
rect -42 36 -36 37
rect -42 29 -41 36
rect -37 29 -36 36
rect -42 28 -36 29
rect -34 36 -28 37
rect -34 29 -33 36
rect -29 29 -28 36
rect -34 28 -28 29
<< ndcontact >>
rect -49 2 -45 6
rect -41 2 -37 6
rect -33 2 -29 6
<< pdcontact >>
rect -49 29 -45 36
rect -41 29 -37 36
rect -33 29 -29 36
<< psubstratepcontact >>
rect -41 -7 -37 -3
<< nsubstratencontact >>
rect -41 41 -37 45
<< polysilicon >>
rect -44 37 -42 39
rect -36 37 -34 39
rect -44 20 -42 28
rect -44 7 -42 16
rect -36 13 -34 28
rect -36 7 -34 9
rect -44 -1 -42 1
rect -36 -1 -34 1
<< polycontact >>
rect -46 16 -42 20
rect -38 9 -34 13
<< metal1 >>
rect -50 41 -41 45
rect -37 41 -28 45
rect -41 36 -37 41
rect -29 29 -28 36
rect -49 26 -46 29
rect -31 26 -28 29
rect -49 23 -28 26
rect -50 16 -46 20
rect -50 9 -38 13
rect -31 6 -28 23
rect -29 2 -28 6
rect -49 -3 -45 2
rect -50 -7 -41 -3
rect -37 -7 -28 -3
<< labels >>
rlabel metal1 -47 43 -47 43 5 vdd
rlabel metal1 -47 -5 -47 -5 1 gnd
rlabel metal1 -29 15 -29 15 1 y
rlabel metal1 -48 18 -48 18 1 a
rlabel metal1 -48 11 -48 11 1 b
<< end >>
