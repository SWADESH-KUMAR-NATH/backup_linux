magic
tech scmos
timestamp 1636469439
<< ntransistor >>
rect -128 -96 -126 -78
rect -120 -96 -118 -78
<< ndiffusion >>
rect -134 -79 -128 -78
rect -134 -95 -133 -79
rect -129 -95 -128 -79
rect -134 -96 -128 -95
rect -126 -79 -120 -78
rect -126 -95 -125 -79
rect -121 -95 -120 -79
rect -126 -96 -120 -95
rect -118 -79 -112 -78
rect -118 -95 -117 -79
rect -113 -95 -112 -79
rect -118 -96 -112 -95
<< ndcontact >>
rect -133 -95 -129 -79
rect -125 -95 -121 -79
rect -117 -95 -113 -79
<< psubstratepcontact >>
rect -125 -74 -121 -70
<< polysilicon >>
rect -128 -78 -126 -76
rect -120 -78 -118 -76
rect -128 -98 -126 -96
rect -120 -98 -118 -96
<< polycontact >>
rect -129 -102 -125 -98
rect -121 -102 -117 -98
<< metal1 >>
rect -148 -74 -125 -70
rect -121 -74 -97 -70
rect -125 -79 -121 -74
rect -136 -85 -133 -81
rect -113 -85 -110 -81
rect -148 -109 -97 -105
rect -136 -134 -122 -130
rect -148 -150 -97 -146
rect -123 -166 -109 -162
rect -148 -191 -97 -187
rect -148 -220 -97 -216
<< m2contact >>
rect -140 -85 -136 -81
rect -110 -85 -106 -81
rect -129 -102 -125 -98
rect -121 -102 -117 -98
rect -141 -118 -137 -114
rect -118 -134 -114 -130
rect -110 -134 -106 -130
rect -108 -158 -104 -154
rect -139 -166 -135 -162
rect -131 -166 -127 -162
rect -121 -206 -117 -202
rect -113 -212 -109 -208
<< metal2 >>
rect -141 -81 -138 -70
rect -108 -81 -105 -70
rect -141 -85 -140 -81
rect -106 -85 -105 -81
rect -128 -115 -125 -102
rect -137 -118 -125 -115
rect -121 -124 -118 -102
rect -121 -127 -100 -124
rect -131 -138 -114 -134
rect -131 -155 -127 -138
rect -110 -141 -106 -134
rect -139 -159 -127 -155
rect -118 -145 -106 -141
rect -139 -162 -135 -159
rect -139 -220 -135 -166
rect -131 -202 -127 -166
rect -118 -167 -114 -145
rect -103 -148 -100 -127
rect -107 -151 -100 -148
rect -107 -154 -104 -151
rect -118 -171 -109 -167
rect -131 -206 -121 -202
rect -131 -220 -127 -206
rect -113 -208 -109 -171
use nand  nand_1
timestamp 1636351123
transform -1 0 -114 0 1 -122
box -17 -28 17 20
use inv  inv_2
timestamp 1636288754
transform -1 0 -135 0 1 -125
box -13 -25 13 23
use nand  nand_2
timestamp 1636351123
transform 1 0 -131 0 -1 -174
box -17 -28 17 20
use inv  inv_1
timestamp 1636288754
transform 1 0 -110 0 -1 -171
box -13 -25 13 23
use inv1  inv1_0
timestamp 1636467228
transform 1 0 -88 0 1 -169
box -48 -51 -9 -15
<< labels >>
rlabel psubstratepcontact -123 -72 -123 -72 1 gnd
rlabel metal2 -140 -77 -140 -77 1 bl
rlabel metal2 -107 -77 -107 -77 1 blb
rlabel metal2 -137 -208 -137 -208 1 w_en
rlabel metal2 -129 -215 -129 -215 1 din
<< end >>
