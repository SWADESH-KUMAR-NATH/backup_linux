magic
tech scmos
timestamp 1636470790
<< nwell >>
rect -257 -57 -215 -19
<< ptransistor >>
rect -245 -43 -243 -25
rect -237 -43 -235 -25
rect -229 -43 -227 -25
<< pdiffusion >>
rect -250 -26 -245 -25
rect -246 -42 -245 -26
rect -250 -43 -245 -42
rect -243 -26 -237 -25
rect -243 -42 -242 -26
rect -238 -42 -237 -26
rect -243 -43 -237 -42
rect -235 -26 -229 -25
rect -235 -42 -234 -26
rect -230 -42 -229 -26
rect -235 -43 -229 -42
rect -227 -26 -222 -25
rect -227 -42 -226 -26
rect -227 -43 -222 -42
<< pdcontact >>
rect -250 -42 -246 -26
rect -242 -42 -238 -26
rect -234 -42 -230 -26
rect -226 -42 -222 -26
<< psubstratepcontact >>
rect -246 -16 -242 -12
rect -230 -16 -226 -12
<< nsubstratencontact >>
rect -246 -54 -242 -50
rect -230 -54 -226 -50
<< polysilicon >>
rect -245 -22 -238 -20
rect -245 -25 -243 -22
rect -234 -22 -227 -20
rect -237 -25 -235 -23
rect -229 -25 -227 -22
rect -245 -45 -243 -43
rect -237 -45 -235 -43
rect -229 -45 -227 -43
<< polycontact >>
rect -238 -23 -234 -19
<< metal1 >>
rect -257 -16 -246 -12
rect -242 -16 -230 -12
rect -226 -16 -215 -12
rect -257 -23 -238 -19
rect -234 -23 -215 -19
rect -250 -50 -246 -42
rect -242 -43 -238 -42
rect -234 -43 -230 -42
rect -226 -50 -222 -42
rect -257 -54 -246 -50
rect -242 -54 -230 -50
rect -226 -54 -215 -50
<< m2contact >>
rect -242 -47 -238 -43
rect -234 -47 -230 -43
<< metal2 >>
rect -254 -47 -242 -43
rect -230 -47 -218 -43
rect -254 -54 -251 -47
rect -221 -54 -218 -47
<< labels >>
rlabel metal1 -236 -52 -236 -52 1 vdd
rlabel metal1 -236 -13 -236 -13 5 gnd
rlabel metal2 -253 -47 -253 -47 3 bl
rlabel metal2 -220 -47 -220 -47 1 blb
rlabel polycontact -236 -21 -236 -21 1 pc
<< end >>
