magic
tech scmos
timestamp 1635858666
<< nwell >>
rect -76 -53 -18 -21
rect -7 -53 61 -12
rect 68 -53 126 -14
<< ptransistor >>
rect -1 -26 17 -24
rect 37 -26 55 -24
rect -56 -45 -54 -27
rect -48 -45 -46 -27
rect -40 -45 -38 -27
rect 26 -47 28 -29
rect 156 -30 165 -28
rect 172 -30 181 -28
rect 188 -30 197 -28
rect 76 -33 85 -31
rect 93 -33 102 -31
rect 109 -33 118 -31
rect 156 -38 165 -36
rect 172 -38 181 -36
rect 188 -38 197 -36
rect 76 -41 85 -39
rect 93 -41 102 -39
rect 109 -41 118 -39
<< pdiffusion >>
rect -1 -19 17 -18
rect -1 -23 0 -19
rect 16 -23 17 -19
rect 37 -19 55 -18
rect 37 -23 38 -19
rect 54 -23 55 -19
rect -1 -24 17 -23
rect -1 -27 17 -26
rect 37 -24 55 -23
rect 156 -23 165 -22
rect 76 -26 85 -25
rect 93 -26 102 -25
rect 37 -27 55 -26
rect -57 -45 -56 -27
rect -54 -45 -53 -27
rect -49 -45 -48 -27
rect -46 -45 -45 -27
rect -41 -45 -40 -27
rect -38 -45 -37 -27
rect -1 -31 0 -27
rect 16 -31 17 -27
rect -1 -32 17 -31
rect 20 -30 26 -29
rect 20 -46 21 -30
rect 25 -46 26 -30
rect 20 -47 26 -46
rect 28 -30 34 -29
rect 28 -46 29 -30
rect 33 -46 34 -30
rect 37 -31 38 -27
rect 54 -31 55 -27
rect 76 -30 77 -26
rect 84 -30 85 -26
rect 76 -31 85 -30
rect 93 -30 94 -26
rect 101 -30 102 -26
rect 93 -31 102 -30
rect 109 -26 118 -25
rect 109 -30 110 -26
rect 117 -30 118 -26
rect 156 -27 157 -23
rect 164 -27 165 -23
rect 156 -28 165 -27
rect 172 -23 181 -22
rect 172 -27 173 -23
rect 180 -27 181 -23
rect 172 -28 181 -27
rect 188 -23 197 -22
rect 188 -27 189 -23
rect 196 -27 197 -23
rect 188 -28 197 -27
rect 109 -31 118 -30
rect 156 -31 165 -30
rect 37 -32 55 -31
rect 76 -34 85 -33
rect 76 -38 77 -34
rect 84 -38 85 -34
rect 76 -39 85 -38
rect 93 -34 102 -33
rect 93 -38 94 -34
rect 101 -38 102 -34
rect 93 -39 102 -38
rect 109 -34 118 -33
rect 109 -38 110 -34
rect 117 -38 118 -34
rect 156 -35 157 -31
rect 164 -35 165 -31
rect 156 -36 165 -35
rect 172 -31 181 -30
rect 172 -35 173 -31
rect 180 -35 181 -31
rect 172 -36 181 -35
rect 188 -31 197 -30
rect 188 -35 189 -31
rect 196 -35 197 -31
rect 188 -36 197 -35
rect 109 -39 118 -38
rect 156 -39 165 -38
rect 28 -47 34 -46
rect 76 -42 85 -41
rect 76 -46 77 -42
rect 84 -46 85 -42
rect 76 -47 85 -46
rect 93 -42 102 -41
rect 93 -46 94 -42
rect 101 -46 102 -42
rect 93 -47 102 -46
rect 109 -42 118 -41
rect 109 -46 110 -42
rect 117 -46 118 -42
rect 156 -43 157 -39
rect 164 -43 165 -39
rect 156 -44 165 -43
rect 172 -39 181 -38
rect 172 -43 173 -39
rect 180 -43 181 -39
rect 172 -44 181 -43
rect 188 -39 197 -38
rect 188 -43 189 -39
rect 196 -43 197 -39
rect 188 -44 197 -43
rect 109 -47 118 -46
<< pdcontact >>
rect 0 -23 16 -19
rect 38 -23 54 -19
rect -61 -45 -57 -27
rect -53 -45 -49 -27
rect -45 -45 -41 -27
rect -37 -45 -33 -27
rect 0 -31 16 -27
rect 21 -46 25 -30
rect 29 -46 33 -30
rect 38 -31 54 -27
rect 77 -30 84 -26
rect 94 -30 101 -26
rect 110 -30 117 -26
rect 157 -27 164 -23
rect 173 -27 180 -23
rect 189 -27 196 -23
rect 77 -38 84 -34
rect 94 -38 101 -34
rect 110 -38 117 -34
rect 157 -35 164 -31
rect 173 -35 180 -31
rect 189 -35 196 -31
rect 77 -46 84 -42
rect 94 -46 101 -42
rect 110 -46 117 -42
rect 157 -43 164 -39
rect 173 -43 180 -39
rect 189 -43 196 -39
<< psubstratepcontact >>
rect 7 -9 11 -5
rect 39 -9 43 -5
rect 79 -11 83 -7
rect 111 -11 115 -7
rect -65 -18 -61 -14
rect -33 -18 -29 -14
<< nsubstratencontact >>
rect 21 -20 25 -16
rect 29 -20 33 -16
rect 72 -21 76 -17
rect 118 -21 122 -17
rect -69 -31 -65 -27
rect -29 -31 -25 -27
<< polysilicon >>
rect -56 -27 -54 -24
rect -48 -27 -46 -24
rect -40 -27 -38 -24
rect -3 -26 -1 -24
rect 17 -26 25 -24
rect 29 -26 37 -24
rect 55 -26 57 -24
rect 26 -29 28 -27
rect -56 -47 -54 -45
rect -48 -47 -46 -45
rect -40 -47 -38 -45
rect 87 -31 91 -30
rect 154 -30 156 -28
rect 165 -30 172 -28
rect 181 -30 188 -28
rect 197 -30 199 -28
rect 74 -33 76 -31
rect 85 -33 93 -31
rect 102 -33 109 -31
rect 118 -33 120 -31
rect 88 -39 90 -33
rect 104 -39 106 -33
rect 154 -38 156 -36
rect 165 -38 172 -36
rect 181 -38 188 -36
rect 197 -38 199 -36
rect 74 -41 76 -39
rect 85 -41 93 -39
rect 102 -41 109 -39
rect 118 -41 120 -39
rect 26 -49 28 -47
<< polycontact >>
rect -57 -24 -53 -20
rect -49 -24 -45 -20
rect -41 -24 -37 -20
rect 25 -27 29 -23
rect 87 -30 91 -26
<< metal1 >>
rect 11 -8 39 -5
rect 83 -10 111 -7
rect -61 -17 -33 -14
rect 0 -19 21 -16
rect -53 -24 -49 -20
rect -45 -24 -41 -20
rect 16 -20 21 -19
rect 25 -20 29 -16
rect 33 -19 54 -16
rect 33 -20 38 -19
rect 71 -21 72 -17
rect 76 -21 80 -17
rect 114 -21 118 -17
rect 122 -21 123 -17
rect 71 -26 74 -21
rect 120 -26 123 -21
rect -65 -30 -61 -27
rect -73 -49 -72 -45
rect -73 -56 -70 -49
rect -61 -52 -57 -45
rect -33 -30 -29 -27
rect 1 -39 4 -31
rect 1 -42 21 -39
rect -37 -52 -33 -45
rect -22 -49 -21 -45
rect -61 -56 -33 -52
rect -24 -56 -21 -49
rect 1 -51 4 -42
rect 71 -30 77 -26
rect 101 -30 107 -26
rect 117 -30 123 -26
rect 50 -39 53 -31
rect 33 -42 53 -39
rect 50 -51 53 -42
rect 71 -42 74 -30
rect 104 -34 107 -30
rect 84 -38 94 -34
rect 104 -38 110 -34
rect 71 -46 77 -42
rect 88 -49 91 -38
rect 104 -42 107 -38
rect 120 -42 123 -30
rect 154 -35 157 -31
rect 101 -46 107 -42
rect 117 -46 123 -42
rect 167 -43 170 -23
rect 183 -43 186 -23
rect 71 -52 91 -49
rect 104 -49 107 -46
rect 104 -52 123 -49
rect 71 -53 74 -52
rect 120 -53 123 -52
<< m2contact >>
rect -57 -24 -53 -20
rect -49 -24 -45 -20
rect -41 -24 -37 -20
rect 80 -21 84 -17
rect 110 -21 114 -17
rect 25 -27 29 -23
rect -72 -49 -68 -45
rect -53 -49 -49 -45
rect -45 -49 -41 -45
rect -26 -49 -22 -45
rect 87 -30 91 -26
<< metal2 >>
rect -76 -17 -18 -14
rect -76 -24 -57 -20
rect -53 -24 -49 -20
rect -45 -24 -41 -20
rect -37 -24 -18 -20
rect 68 -21 80 -17
rect 84 -21 110 -17
rect 114 -21 126 -17
rect -7 -27 25 -23
rect 29 -27 61 -23
rect 68 -30 87 -26
rect 91 -30 126 -26
rect -68 -49 -53 -45
rect -41 -49 -26 -45
rect -76 -56 -18 -52
use pc  pc_0
timestamp 1635740445
transform 1 0 -171 0 1 -4
box 0 -47 58 -8
<< labels >>
rlabel metal1 -23 -50 -22 -49 8 blb
rlabel metal1 -72 -50 -71 -49 2 bl
rlabel metal1 -47 -15 -47 -15 5 gnd
rlabel metal1 25 -6 25 -6 5 gnd
rlabel metal1 97 -8 97 -8 5 gnd
rlabel metal2 -73 -22 -73 -22 3 pc
rlabel metal1 -47 -54 -47 -54 1 vdd
<< end >>
