magic
tech scmos
timestamp 1636470524
<< nwell >>
rect -191 27 -149 48
<< ntransistor >>
rect -175 13 -173 19
rect -167 13 -165 19
rect -179 4 -176 8
rect -164 4 -161 8
<< ptransistor >>
rect -179 34 -173 37
rect -167 34 -161 37
<< ndiffusion >>
rect -181 18 -175 19
rect -181 14 -180 18
rect -176 14 -175 18
rect -181 13 -175 14
rect -173 18 -167 19
rect -173 14 -172 18
rect -168 14 -167 18
rect -173 13 -167 14
rect -165 18 -159 19
rect -165 14 -164 18
rect -160 14 -159 18
rect -165 13 -159 14
rect -179 8 -176 13
rect -164 8 -161 13
rect -179 3 -176 4
rect -164 3 -161 4
<< pdiffusion >>
rect -180 34 -179 37
rect -173 35 -172 37
rect -168 35 -167 37
rect -173 34 -167 35
rect -161 34 -160 37
<< ndcontact >>
rect -180 14 -176 18
rect -172 14 -168 18
rect -164 14 -160 18
rect -180 -1 -176 3
rect -164 -1 -160 3
<< pdcontact >>
rect -184 33 -180 37
rect -172 35 -168 39
rect -160 33 -156 37
<< psubstratepcontact >>
rect -172 -8 -168 -4
<< nsubstratencontact >>
rect -180 41 -176 45
rect -164 41 -160 45
<< polysilicon >>
rect -179 37 -173 39
rect -167 37 -161 39
rect -179 32 -173 34
rect -167 32 -161 34
rect -175 19 -173 28
rect -167 25 -165 32
rect -167 19 -165 21
rect -175 11 -173 13
rect -167 11 -165 13
rect -180 6 -179 8
rect -184 4 -179 6
rect -176 4 -164 8
rect -161 6 -160 8
rect -161 4 -156 6
<< polycontact >>
rect -175 28 -171 32
rect -169 21 -165 25
rect -184 6 -180 10
rect -160 6 -156 10
<< metal1 >>
rect -191 41 -180 45
rect -176 41 -164 45
rect -160 41 -149 45
rect -172 39 -168 41
rect -183 31 -180 33
rect -183 28 -178 31
rect -160 31 -157 33
rect -171 28 -157 31
rect -181 25 -178 28
rect -181 22 -169 25
rect -181 18 -178 22
rect -162 18 -159 28
rect -181 14 -180 18
rect -160 14 -159 18
rect -191 6 -184 10
rect -181 -1 -180 3
rect -172 -4 -168 14
rect -156 6 -149 10
rect -160 -1 -159 3
rect -191 -8 -172 -4
rect -168 -8 -149 -4
<< m2contact >>
rect -185 -1 -181 3
rect -159 -1 -155 3
<< metal2 >>
rect -188 -8 -185 48
rect -155 -8 -152 48
<< labels >>
rlabel metal1 -170 43 -170 43 5 vdd
rlabel psubstratepcontact -170 -6 -170 -6 1 gnd
rlabel metal1 -189 8 -189 8 3 wl
rlabel metal2 -187 20 -187 20 3 bl
rlabel metal2 -153 20 -153 20 7 blb
rlabel metal1 -179 23 -179 23 1 q1
rlabel metal1 -161 23 -161 23 1 q2
<< end >>
