magic
tech scmos
timestamp 1633895608
<< nwell >>
rect -13 -4 13 23
<< ntransistor >>
rect -1 -14 1 -10
<< ptransistor >>
rect -1 2 1 12
<< ndiffusion >>
rect -7 -14 -6 -10
rect -2 -14 -1 -10
rect 1 -14 2 -10
rect 6 -14 7 -10
<< pdiffusion >>
rect -7 11 -1 12
rect -7 3 -6 11
rect -2 3 -1 11
rect -7 2 -1 3
rect 1 11 7 12
rect 1 3 2 11
rect 6 3 7 11
rect 1 2 7 3
<< ndcontact >>
rect -6 -14 -2 -10
rect 2 -14 6 -10
<< pdcontact >>
rect -6 3 -2 11
rect 2 3 6 11
<< psubstratepcontact >>
rect -6 -22 -2 -18
rect 2 -22 6 -18
<< nsubstratencontact >>
rect -6 16 -2 20
rect 2 16 6 20
<< polysilicon >>
rect -1 12 1 14
rect -1 -2 1 2
rect 0 -6 1 -2
rect -1 -10 1 -6
rect -1 -16 1 -14
<< polycontact >>
rect -4 -6 0 -2
<< metal1 >>
rect -7 16 -6 20
rect -2 16 2 20
rect 6 16 7 20
rect -6 11 -2 16
rect -7 -6 -4 -2
rect 3 -10 6 3
rect -6 -18 -2 -14
rect -7 -22 -6 -18
rect -2 -22 2 -18
rect 6 -22 7 -18
<< labels >>
rlabel metal1 -6 -4 -6 -4 1 in
rlabel metal1 4 -4 4 -4 1 out
<< end >>
