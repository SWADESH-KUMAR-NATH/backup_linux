magic
tech scmos
timestamp 1635858666
<< nwell >>
rect 198 -110 641 -89
rect 198 -182 641 -150
rect 198 -254 641 -222
rect 198 -326 641 -294
rect 198 -387 641 -366
<< ntransistor >>
rect 207 -122 211 -119
rect 222 -124 224 -118
rect 230 -124 232 -118
rect 243 -122 247 -119
rect 262 -122 266 -119
rect 277 -124 279 -118
rect 285 -124 287 -118
rect 298 -122 302 -119
rect 317 -122 321 -119
rect 332 -124 334 -118
rect 340 -124 342 -118
rect 353 -122 357 -119
rect 372 -122 376 -119
rect 387 -124 389 -118
rect 395 -124 397 -118
rect 408 -122 412 -119
rect 427 -122 431 -119
rect 442 -124 444 -118
rect 450 -124 452 -118
rect 463 -122 467 -119
rect 482 -122 486 -119
rect 497 -124 499 -118
rect 505 -124 507 -118
rect 518 -122 522 -119
rect 537 -122 541 -119
rect 552 -124 554 -118
rect 560 -124 562 -118
rect 573 -122 577 -119
rect 592 -122 596 -119
rect 607 -124 609 -118
rect 615 -124 617 -118
rect 628 -122 632 -119
rect 207 -141 211 -138
rect 222 -142 224 -136
rect 230 -142 232 -136
rect 243 -141 247 -138
rect 262 -141 266 -138
rect 277 -142 279 -136
rect 285 -142 287 -136
rect 298 -141 302 -138
rect 317 -141 321 -138
rect 332 -142 334 -136
rect 340 -142 342 -136
rect 353 -141 357 -138
rect 372 -141 376 -138
rect 387 -142 389 -136
rect 395 -142 397 -136
rect 408 -141 412 -138
rect 427 -141 431 -138
rect 442 -142 444 -136
rect 450 -142 452 -136
rect 463 -141 467 -138
rect 482 -141 486 -138
rect 497 -142 499 -136
rect 505 -142 507 -136
rect 518 -141 522 -138
rect 537 -141 541 -138
rect 552 -142 554 -136
rect 560 -142 562 -136
rect 573 -141 577 -138
rect 592 -141 596 -138
rect 607 -142 609 -136
rect 615 -142 617 -136
rect 628 -141 632 -138
rect 207 -194 211 -191
rect 222 -196 224 -190
rect 230 -196 232 -190
rect 243 -194 247 -191
rect 262 -194 266 -191
rect 277 -196 279 -190
rect 285 -196 287 -190
rect 298 -194 302 -191
rect 317 -194 321 -191
rect 332 -196 334 -190
rect 340 -196 342 -190
rect 353 -194 357 -191
rect 372 -194 376 -191
rect 387 -196 389 -190
rect 395 -196 397 -190
rect 408 -194 412 -191
rect 427 -194 431 -191
rect 442 -196 444 -190
rect 450 -196 452 -190
rect 463 -194 467 -191
rect 482 -194 486 -191
rect 497 -196 499 -190
rect 505 -196 507 -190
rect 518 -194 522 -191
rect 537 -194 541 -191
rect 552 -196 554 -190
rect 560 -196 562 -190
rect 573 -194 577 -191
rect 592 -194 596 -191
rect 607 -196 609 -190
rect 615 -196 617 -190
rect 628 -194 632 -191
rect 207 -213 211 -210
rect 222 -214 224 -208
rect 230 -214 232 -208
rect 243 -213 247 -210
rect 262 -213 266 -210
rect 277 -214 279 -208
rect 285 -214 287 -208
rect 298 -213 302 -210
rect 317 -213 321 -210
rect 332 -214 334 -208
rect 340 -214 342 -208
rect 353 -213 357 -210
rect 372 -213 376 -210
rect 387 -214 389 -208
rect 395 -214 397 -208
rect 408 -213 412 -210
rect 427 -213 431 -210
rect 442 -214 444 -208
rect 450 -214 452 -208
rect 463 -213 467 -210
rect 482 -213 486 -210
rect 497 -214 499 -208
rect 505 -214 507 -208
rect 518 -213 522 -210
rect 537 -213 541 -210
rect 552 -214 554 -208
rect 560 -214 562 -208
rect 573 -213 577 -210
rect 592 -213 596 -210
rect 607 -214 609 -208
rect 615 -214 617 -208
rect 628 -213 632 -210
rect 207 -266 211 -263
rect 222 -268 224 -262
rect 230 -268 232 -262
rect 243 -266 247 -263
rect 262 -266 266 -263
rect 277 -268 279 -262
rect 285 -268 287 -262
rect 298 -266 302 -263
rect 317 -266 321 -263
rect 332 -268 334 -262
rect 340 -268 342 -262
rect 353 -266 357 -263
rect 372 -266 376 -263
rect 387 -268 389 -262
rect 395 -268 397 -262
rect 408 -266 412 -263
rect 427 -266 431 -263
rect 442 -268 444 -262
rect 450 -268 452 -262
rect 463 -266 467 -263
rect 482 -266 486 -263
rect 497 -268 499 -262
rect 505 -268 507 -262
rect 518 -266 522 -263
rect 537 -266 541 -263
rect 552 -268 554 -262
rect 560 -268 562 -262
rect 573 -266 577 -263
rect 592 -266 596 -263
rect 607 -268 609 -262
rect 615 -268 617 -262
rect 628 -266 632 -263
rect 207 -285 211 -282
rect 222 -286 224 -280
rect 230 -286 232 -280
rect 243 -285 247 -282
rect 262 -285 266 -282
rect 277 -286 279 -280
rect 285 -286 287 -280
rect 298 -285 302 -282
rect 317 -285 321 -282
rect 332 -286 334 -280
rect 340 -286 342 -280
rect 353 -285 357 -282
rect 372 -285 376 -282
rect 387 -286 389 -280
rect 395 -286 397 -280
rect 408 -285 412 -282
rect 427 -285 431 -282
rect 442 -286 444 -280
rect 450 -286 452 -280
rect 463 -285 467 -282
rect 482 -285 486 -282
rect 497 -286 499 -280
rect 505 -286 507 -280
rect 518 -285 522 -282
rect 537 -285 541 -282
rect 552 -286 554 -280
rect 560 -286 562 -280
rect 573 -285 577 -282
rect 592 -285 596 -282
rect 607 -286 609 -280
rect 615 -286 617 -280
rect 628 -285 632 -282
rect 207 -338 211 -335
rect 222 -340 224 -334
rect 230 -340 232 -334
rect 243 -338 247 -335
rect 262 -338 266 -335
rect 277 -340 279 -334
rect 285 -340 287 -334
rect 298 -338 302 -335
rect 317 -338 321 -335
rect 332 -340 334 -334
rect 340 -340 342 -334
rect 353 -338 357 -335
rect 372 -338 376 -335
rect 387 -340 389 -334
rect 395 -340 397 -334
rect 408 -338 412 -335
rect 427 -338 431 -335
rect 442 -340 444 -334
rect 450 -340 452 -334
rect 463 -338 467 -335
rect 482 -338 486 -335
rect 497 -340 499 -334
rect 505 -340 507 -334
rect 518 -338 522 -335
rect 537 -338 541 -335
rect 552 -340 554 -334
rect 560 -340 562 -334
rect 573 -338 577 -335
rect 592 -338 596 -335
rect 607 -340 609 -334
rect 615 -340 617 -334
rect 628 -338 632 -335
rect 207 -357 211 -354
rect 222 -358 224 -352
rect 230 -358 232 -352
rect 243 -357 247 -354
rect 262 -357 266 -354
rect 277 -358 279 -352
rect 285 -358 287 -352
rect 298 -357 302 -354
rect 317 -357 321 -354
rect 332 -358 334 -352
rect 340 -358 342 -352
rect 353 -357 357 -354
rect 372 -357 376 -354
rect 387 -358 389 -352
rect 395 -358 397 -352
rect 408 -357 412 -354
rect 427 -357 431 -354
rect 442 -358 444 -352
rect 450 -358 452 -352
rect 463 -357 467 -354
rect 482 -357 486 -354
rect 497 -358 499 -352
rect 505 -358 507 -352
rect 518 -357 522 -354
rect 537 -357 541 -354
rect 552 -358 554 -352
rect 560 -358 562 -352
rect 573 -357 577 -354
rect 592 -357 596 -354
rect 607 -358 609 -352
rect 615 -358 617 -352
rect 628 -357 632 -354
<< ptransistor >>
rect 218 -103 224 -100
rect 230 -103 236 -100
rect 273 -103 279 -100
rect 285 -103 291 -100
rect 328 -103 334 -100
rect 340 -103 346 -100
rect 383 -103 389 -100
rect 395 -103 401 -100
rect 438 -103 444 -100
rect 450 -103 456 -100
rect 493 -103 499 -100
rect 505 -103 511 -100
rect 548 -103 554 -100
rect 560 -103 566 -100
rect 603 -103 609 -100
rect 615 -103 621 -100
rect 218 -160 224 -157
rect 230 -160 236 -157
rect 273 -160 279 -157
rect 285 -160 291 -157
rect 328 -160 334 -157
rect 340 -160 346 -157
rect 383 -160 389 -157
rect 395 -160 401 -157
rect 438 -160 444 -157
rect 450 -160 456 -157
rect 493 -160 499 -157
rect 505 -160 511 -157
rect 548 -160 554 -157
rect 560 -160 566 -157
rect 603 -160 609 -157
rect 615 -160 621 -157
rect 218 -175 224 -172
rect 230 -175 236 -172
rect 273 -175 279 -172
rect 285 -175 291 -172
rect 328 -175 334 -172
rect 340 -175 346 -172
rect 383 -175 389 -172
rect 395 -175 401 -172
rect 438 -175 444 -172
rect 450 -175 456 -172
rect 493 -175 499 -172
rect 505 -175 511 -172
rect 548 -175 554 -172
rect 560 -175 566 -172
rect 603 -175 609 -172
rect 615 -175 621 -172
rect 218 -232 224 -229
rect 230 -232 236 -229
rect 273 -232 279 -229
rect 285 -232 291 -229
rect 328 -232 334 -229
rect 340 -232 346 -229
rect 383 -232 389 -229
rect 395 -232 401 -229
rect 438 -232 444 -229
rect 450 -232 456 -229
rect 493 -232 499 -229
rect 505 -232 511 -229
rect 548 -232 554 -229
rect 560 -232 566 -229
rect 603 -232 609 -229
rect 615 -232 621 -229
rect 218 -247 224 -244
rect 230 -247 236 -244
rect 273 -247 279 -244
rect 285 -247 291 -244
rect 328 -247 334 -244
rect 340 -247 346 -244
rect 383 -247 389 -244
rect 395 -247 401 -244
rect 438 -247 444 -244
rect 450 -247 456 -244
rect 493 -247 499 -244
rect 505 -247 511 -244
rect 548 -247 554 -244
rect 560 -247 566 -244
rect 603 -247 609 -244
rect 615 -247 621 -244
rect 218 -304 224 -301
rect 230 -304 236 -301
rect 273 -304 279 -301
rect 285 -304 291 -301
rect 328 -304 334 -301
rect 340 -304 346 -301
rect 383 -304 389 -301
rect 395 -304 401 -301
rect 438 -304 444 -301
rect 450 -304 456 -301
rect 493 -304 499 -301
rect 505 -304 511 -301
rect 548 -304 554 -301
rect 560 -304 566 -301
rect 603 -304 609 -301
rect 615 -304 621 -301
rect 218 -319 224 -316
rect 230 -319 236 -316
rect 273 -319 279 -316
rect 285 -319 291 -316
rect 328 -319 334 -316
rect 340 -319 346 -316
rect 383 -319 389 -316
rect 395 -319 401 -316
rect 438 -319 444 -316
rect 450 -319 456 -316
rect 493 -319 499 -316
rect 505 -319 511 -316
rect 548 -319 554 -316
rect 560 -319 566 -316
rect 603 -319 609 -316
rect 615 -319 621 -316
rect 218 -376 224 -373
rect 230 -376 236 -373
rect 273 -376 279 -373
rect 285 -376 291 -373
rect 328 -376 334 -373
rect 340 -376 346 -373
rect 383 -376 389 -373
rect 395 -376 401 -373
rect 438 -376 444 -373
rect 450 -376 456 -373
rect 493 -376 499 -373
rect 505 -376 511 -373
rect 548 -376 554 -373
rect 560 -376 566 -373
rect 603 -376 609 -373
rect 615 -376 621 -373
<< ndiffusion >>
rect 212 -119 222 -118
rect 206 -122 207 -119
rect 211 -122 212 -119
rect 219 -123 222 -119
rect 212 -124 222 -123
rect 224 -119 230 -118
rect 224 -123 225 -119
rect 229 -123 230 -119
rect 224 -124 230 -123
rect 232 -119 242 -118
rect 267 -119 277 -118
rect 232 -123 235 -119
rect 242 -122 243 -119
rect 247 -122 248 -119
rect 232 -124 242 -123
rect 261 -122 262 -119
rect 266 -122 267 -119
rect 274 -123 277 -119
rect 267 -124 277 -123
rect 279 -119 285 -118
rect 279 -123 280 -119
rect 284 -123 285 -119
rect 279 -124 285 -123
rect 287 -119 297 -118
rect 322 -119 332 -118
rect 287 -123 290 -119
rect 297 -122 298 -119
rect 302 -122 303 -119
rect 287 -124 297 -123
rect 316 -122 317 -119
rect 321 -122 322 -119
rect 329 -123 332 -119
rect 322 -124 332 -123
rect 334 -119 340 -118
rect 334 -123 335 -119
rect 339 -123 340 -119
rect 334 -124 340 -123
rect 342 -119 352 -118
rect 377 -119 387 -118
rect 342 -123 345 -119
rect 352 -122 353 -119
rect 357 -122 358 -119
rect 342 -124 352 -123
rect 371 -122 372 -119
rect 376 -122 377 -119
rect 384 -123 387 -119
rect 377 -124 387 -123
rect 389 -119 395 -118
rect 389 -123 390 -119
rect 394 -123 395 -119
rect 389 -124 395 -123
rect 397 -119 407 -118
rect 432 -119 442 -118
rect 397 -123 400 -119
rect 407 -122 408 -119
rect 412 -122 413 -119
rect 397 -124 407 -123
rect 426 -122 427 -119
rect 431 -122 432 -119
rect 439 -123 442 -119
rect 432 -124 442 -123
rect 444 -119 450 -118
rect 444 -123 445 -119
rect 449 -123 450 -119
rect 444 -124 450 -123
rect 452 -119 462 -118
rect 487 -119 497 -118
rect 452 -123 455 -119
rect 462 -122 463 -119
rect 467 -122 468 -119
rect 452 -124 462 -123
rect 481 -122 482 -119
rect 486 -122 487 -119
rect 494 -123 497 -119
rect 487 -124 497 -123
rect 499 -119 505 -118
rect 499 -123 500 -119
rect 504 -123 505 -119
rect 499 -124 505 -123
rect 507 -119 517 -118
rect 542 -119 552 -118
rect 507 -123 510 -119
rect 517 -122 518 -119
rect 522 -122 523 -119
rect 507 -124 517 -123
rect 536 -122 537 -119
rect 541 -122 542 -119
rect 549 -123 552 -119
rect 542 -124 552 -123
rect 554 -119 560 -118
rect 554 -123 555 -119
rect 559 -123 560 -119
rect 554 -124 560 -123
rect 562 -119 572 -118
rect 597 -119 607 -118
rect 562 -123 565 -119
rect 572 -122 573 -119
rect 577 -122 578 -119
rect 562 -124 572 -123
rect 591 -122 592 -119
rect 596 -122 597 -119
rect 604 -123 607 -119
rect 597 -124 607 -123
rect 609 -119 615 -118
rect 609 -123 610 -119
rect 614 -123 615 -119
rect 609 -124 615 -123
rect 617 -119 627 -118
rect 617 -123 620 -119
rect 627 -122 628 -119
rect 632 -122 633 -119
rect 617 -124 627 -123
rect 212 -137 222 -136
rect 206 -141 207 -138
rect 211 -141 212 -138
rect 219 -141 222 -137
rect 212 -142 222 -141
rect 224 -137 230 -136
rect 224 -141 225 -137
rect 229 -141 230 -137
rect 224 -142 230 -141
rect 232 -137 242 -136
rect 232 -141 235 -137
rect 242 -141 243 -138
rect 247 -141 248 -138
rect 267 -137 277 -136
rect 261 -141 262 -138
rect 266 -141 267 -138
rect 274 -141 277 -137
rect 232 -142 242 -141
rect 267 -142 277 -141
rect 279 -137 285 -136
rect 279 -141 280 -137
rect 284 -141 285 -137
rect 279 -142 285 -141
rect 287 -137 297 -136
rect 287 -141 290 -137
rect 297 -141 298 -138
rect 302 -141 303 -138
rect 322 -137 332 -136
rect 316 -141 317 -138
rect 321 -141 322 -138
rect 329 -141 332 -137
rect 287 -142 297 -141
rect 322 -142 332 -141
rect 334 -137 340 -136
rect 334 -141 335 -137
rect 339 -141 340 -137
rect 334 -142 340 -141
rect 342 -137 352 -136
rect 342 -141 345 -137
rect 352 -141 353 -138
rect 357 -141 358 -138
rect 377 -137 387 -136
rect 371 -141 372 -138
rect 376 -141 377 -138
rect 384 -141 387 -137
rect 342 -142 352 -141
rect 377 -142 387 -141
rect 389 -137 395 -136
rect 389 -141 390 -137
rect 394 -141 395 -137
rect 389 -142 395 -141
rect 397 -137 407 -136
rect 397 -141 400 -137
rect 407 -141 408 -138
rect 412 -141 413 -138
rect 432 -137 442 -136
rect 426 -141 427 -138
rect 431 -141 432 -138
rect 439 -141 442 -137
rect 397 -142 407 -141
rect 432 -142 442 -141
rect 444 -137 450 -136
rect 444 -141 445 -137
rect 449 -141 450 -137
rect 444 -142 450 -141
rect 452 -137 462 -136
rect 452 -141 455 -137
rect 462 -141 463 -138
rect 467 -141 468 -138
rect 487 -137 497 -136
rect 481 -141 482 -138
rect 486 -141 487 -138
rect 494 -141 497 -137
rect 452 -142 462 -141
rect 487 -142 497 -141
rect 499 -137 505 -136
rect 499 -141 500 -137
rect 504 -141 505 -137
rect 499 -142 505 -141
rect 507 -137 517 -136
rect 507 -141 510 -137
rect 517 -141 518 -138
rect 522 -141 523 -138
rect 542 -137 552 -136
rect 536 -141 537 -138
rect 541 -141 542 -138
rect 549 -141 552 -137
rect 507 -142 517 -141
rect 542 -142 552 -141
rect 554 -137 560 -136
rect 554 -141 555 -137
rect 559 -141 560 -137
rect 554 -142 560 -141
rect 562 -137 572 -136
rect 562 -141 565 -137
rect 572 -141 573 -138
rect 577 -141 578 -138
rect 597 -137 607 -136
rect 591 -141 592 -138
rect 596 -141 597 -138
rect 604 -141 607 -137
rect 562 -142 572 -141
rect 597 -142 607 -141
rect 609 -137 615 -136
rect 609 -141 610 -137
rect 614 -141 615 -137
rect 609 -142 615 -141
rect 617 -137 627 -136
rect 617 -141 620 -137
rect 627 -141 628 -138
rect 632 -141 633 -138
rect 617 -142 627 -141
rect 212 -191 222 -190
rect 206 -194 207 -191
rect 211 -194 212 -191
rect 219 -195 222 -191
rect 212 -196 222 -195
rect 224 -191 230 -190
rect 224 -195 225 -191
rect 229 -195 230 -191
rect 224 -196 230 -195
rect 232 -191 242 -190
rect 267 -191 277 -190
rect 232 -195 235 -191
rect 242 -194 243 -191
rect 247 -194 248 -191
rect 232 -196 242 -195
rect 261 -194 262 -191
rect 266 -194 267 -191
rect 274 -195 277 -191
rect 267 -196 277 -195
rect 279 -191 285 -190
rect 279 -195 280 -191
rect 284 -195 285 -191
rect 279 -196 285 -195
rect 287 -191 297 -190
rect 322 -191 332 -190
rect 287 -195 290 -191
rect 297 -194 298 -191
rect 302 -194 303 -191
rect 287 -196 297 -195
rect 316 -194 317 -191
rect 321 -194 322 -191
rect 329 -195 332 -191
rect 322 -196 332 -195
rect 334 -191 340 -190
rect 334 -195 335 -191
rect 339 -195 340 -191
rect 334 -196 340 -195
rect 342 -191 352 -190
rect 377 -191 387 -190
rect 342 -195 345 -191
rect 352 -194 353 -191
rect 357 -194 358 -191
rect 342 -196 352 -195
rect 371 -194 372 -191
rect 376 -194 377 -191
rect 384 -195 387 -191
rect 377 -196 387 -195
rect 389 -191 395 -190
rect 389 -195 390 -191
rect 394 -195 395 -191
rect 389 -196 395 -195
rect 397 -191 407 -190
rect 432 -191 442 -190
rect 397 -195 400 -191
rect 407 -194 408 -191
rect 412 -194 413 -191
rect 397 -196 407 -195
rect 426 -194 427 -191
rect 431 -194 432 -191
rect 439 -195 442 -191
rect 432 -196 442 -195
rect 444 -191 450 -190
rect 444 -195 445 -191
rect 449 -195 450 -191
rect 444 -196 450 -195
rect 452 -191 462 -190
rect 487 -191 497 -190
rect 452 -195 455 -191
rect 462 -194 463 -191
rect 467 -194 468 -191
rect 452 -196 462 -195
rect 481 -194 482 -191
rect 486 -194 487 -191
rect 494 -195 497 -191
rect 487 -196 497 -195
rect 499 -191 505 -190
rect 499 -195 500 -191
rect 504 -195 505 -191
rect 499 -196 505 -195
rect 507 -191 517 -190
rect 542 -191 552 -190
rect 507 -195 510 -191
rect 517 -194 518 -191
rect 522 -194 523 -191
rect 507 -196 517 -195
rect 536 -194 537 -191
rect 541 -194 542 -191
rect 549 -195 552 -191
rect 542 -196 552 -195
rect 554 -191 560 -190
rect 554 -195 555 -191
rect 559 -195 560 -191
rect 554 -196 560 -195
rect 562 -191 572 -190
rect 597 -191 607 -190
rect 562 -195 565 -191
rect 572 -194 573 -191
rect 577 -194 578 -191
rect 562 -196 572 -195
rect 591 -194 592 -191
rect 596 -194 597 -191
rect 604 -195 607 -191
rect 597 -196 607 -195
rect 609 -191 615 -190
rect 609 -195 610 -191
rect 614 -195 615 -191
rect 609 -196 615 -195
rect 617 -191 627 -190
rect 617 -195 620 -191
rect 627 -194 628 -191
rect 632 -194 633 -191
rect 617 -196 627 -195
rect 212 -209 222 -208
rect 206 -213 207 -210
rect 211 -213 212 -210
rect 219 -213 222 -209
rect 212 -214 222 -213
rect 224 -209 230 -208
rect 224 -213 225 -209
rect 229 -213 230 -209
rect 224 -214 230 -213
rect 232 -209 242 -208
rect 232 -213 235 -209
rect 242 -213 243 -210
rect 247 -213 248 -210
rect 267 -209 277 -208
rect 261 -213 262 -210
rect 266 -213 267 -210
rect 274 -213 277 -209
rect 232 -214 242 -213
rect 267 -214 277 -213
rect 279 -209 285 -208
rect 279 -213 280 -209
rect 284 -213 285 -209
rect 279 -214 285 -213
rect 287 -209 297 -208
rect 287 -213 290 -209
rect 297 -213 298 -210
rect 302 -213 303 -210
rect 322 -209 332 -208
rect 316 -213 317 -210
rect 321 -213 322 -210
rect 329 -213 332 -209
rect 287 -214 297 -213
rect 322 -214 332 -213
rect 334 -209 340 -208
rect 334 -213 335 -209
rect 339 -213 340 -209
rect 334 -214 340 -213
rect 342 -209 352 -208
rect 342 -213 345 -209
rect 352 -213 353 -210
rect 357 -213 358 -210
rect 377 -209 387 -208
rect 371 -213 372 -210
rect 376 -213 377 -210
rect 384 -213 387 -209
rect 342 -214 352 -213
rect 377 -214 387 -213
rect 389 -209 395 -208
rect 389 -213 390 -209
rect 394 -213 395 -209
rect 389 -214 395 -213
rect 397 -209 407 -208
rect 397 -213 400 -209
rect 407 -213 408 -210
rect 412 -213 413 -210
rect 432 -209 442 -208
rect 426 -213 427 -210
rect 431 -213 432 -210
rect 439 -213 442 -209
rect 397 -214 407 -213
rect 432 -214 442 -213
rect 444 -209 450 -208
rect 444 -213 445 -209
rect 449 -213 450 -209
rect 444 -214 450 -213
rect 452 -209 462 -208
rect 452 -213 455 -209
rect 462 -213 463 -210
rect 467 -213 468 -210
rect 487 -209 497 -208
rect 481 -213 482 -210
rect 486 -213 487 -210
rect 494 -213 497 -209
rect 452 -214 462 -213
rect 487 -214 497 -213
rect 499 -209 505 -208
rect 499 -213 500 -209
rect 504 -213 505 -209
rect 499 -214 505 -213
rect 507 -209 517 -208
rect 507 -213 510 -209
rect 517 -213 518 -210
rect 522 -213 523 -210
rect 542 -209 552 -208
rect 536 -213 537 -210
rect 541 -213 542 -210
rect 549 -213 552 -209
rect 507 -214 517 -213
rect 542 -214 552 -213
rect 554 -209 560 -208
rect 554 -213 555 -209
rect 559 -213 560 -209
rect 554 -214 560 -213
rect 562 -209 572 -208
rect 562 -213 565 -209
rect 572 -213 573 -210
rect 577 -213 578 -210
rect 597 -209 607 -208
rect 591 -213 592 -210
rect 596 -213 597 -210
rect 604 -213 607 -209
rect 562 -214 572 -213
rect 597 -214 607 -213
rect 609 -209 615 -208
rect 609 -213 610 -209
rect 614 -213 615 -209
rect 609 -214 615 -213
rect 617 -209 627 -208
rect 617 -213 620 -209
rect 627 -213 628 -210
rect 632 -213 633 -210
rect 617 -214 627 -213
rect 212 -263 222 -262
rect 206 -266 207 -263
rect 211 -266 212 -263
rect 219 -267 222 -263
rect 212 -268 222 -267
rect 224 -263 230 -262
rect 224 -267 225 -263
rect 229 -267 230 -263
rect 224 -268 230 -267
rect 232 -263 242 -262
rect 267 -263 277 -262
rect 232 -267 235 -263
rect 242 -266 243 -263
rect 247 -266 248 -263
rect 232 -268 242 -267
rect 261 -266 262 -263
rect 266 -266 267 -263
rect 274 -267 277 -263
rect 267 -268 277 -267
rect 279 -263 285 -262
rect 279 -267 280 -263
rect 284 -267 285 -263
rect 279 -268 285 -267
rect 287 -263 297 -262
rect 322 -263 332 -262
rect 287 -267 290 -263
rect 297 -266 298 -263
rect 302 -266 303 -263
rect 287 -268 297 -267
rect 316 -266 317 -263
rect 321 -266 322 -263
rect 329 -267 332 -263
rect 322 -268 332 -267
rect 334 -263 340 -262
rect 334 -267 335 -263
rect 339 -267 340 -263
rect 334 -268 340 -267
rect 342 -263 352 -262
rect 377 -263 387 -262
rect 342 -267 345 -263
rect 352 -266 353 -263
rect 357 -266 358 -263
rect 342 -268 352 -267
rect 371 -266 372 -263
rect 376 -266 377 -263
rect 384 -267 387 -263
rect 377 -268 387 -267
rect 389 -263 395 -262
rect 389 -267 390 -263
rect 394 -267 395 -263
rect 389 -268 395 -267
rect 397 -263 407 -262
rect 432 -263 442 -262
rect 397 -267 400 -263
rect 407 -266 408 -263
rect 412 -266 413 -263
rect 397 -268 407 -267
rect 426 -266 427 -263
rect 431 -266 432 -263
rect 439 -267 442 -263
rect 432 -268 442 -267
rect 444 -263 450 -262
rect 444 -267 445 -263
rect 449 -267 450 -263
rect 444 -268 450 -267
rect 452 -263 462 -262
rect 487 -263 497 -262
rect 452 -267 455 -263
rect 462 -266 463 -263
rect 467 -266 468 -263
rect 452 -268 462 -267
rect 481 -266 482 -263
rect 486 -266 487 -263
rect 494 -267 497 -263
rect 487 -268 497 -267
rect 499 -263 505 -262
rect 499 -267 500 -263
rect 504 -267 505 -263
rect 499 -268 505 -267
rect 507 -263 517 -262
rect 542 -263 552 -262
rect 507 -267 510 -263
rect 517 -266 518 -263
rect 522 -266 523 -263
rect 507 -268 517 -267
rect 536 -266 537 -263
rect 541 -266 542 -263
rect 549 -267 552 -263
rect 542 -268 552 -267
rect 554 -263 560 -262
rect 554 -267 555 -263
rect 559 -267 560 -263
rect 554 -268 560 -267
rect 562 -263 572 -262
rect 597 -263 607 -262
rect 562 -267 565 -263
rect 572 -266 573 -263
rect 577 -266 578 -263
rect 562 -268 572 -267
rect 591 -266 592 -263
rect 596 -266 597 -263
rect 604 -267 607 -263
rect 597 -268 607 -267
rect 609 -263 615 -262
rect 609 -267 610 -263
rect 614 -267 615 -263
rect 609 -268 615 -267
rect 617 -263 627 -262
rect 617 -267 620 -263
rect 627 -266 628 -263
rect 632 -266 633 -263
rect 617 -268 627 -267
rect 212 -281 222 -280
rect 206 -285 207 -282
rect 211 -285 212 -282
rect 219 -285 222 -281
rect 212 -286 222 -285
rect 224 -281 230 -280
rect 224 -285 225 -281
rect 229 -285 230 -281
rect 224 -286 230 -285
rect 232 -281 242 -280
rect 232 -285 235 -281
rect 242 -285 243 -282
rect 247 -285 248 -282
rect 267 -281 277 -280
rect 261 -285 262 -282
rect 266 -285 267 -282
rect 274 -285 277 -281
rect 232 -286 242 -285
rect 267 -286 277 -285
rect 279 -281 285 -280
rect 279 -285 280 -281
rect 284 -285 285 -281
rect 279 -286 285 -285
rect 287 -281 297 -280
rect 287 -285 290 -281
rect 297 -285 298 -282
rect 302 -285 303 -282
rect 322 -281 332 -280
rect 316 -285 317 -282
rect 321 -285 322 -282
rect 329 -285 332 -281
rect 287 -286 297 -285
rect 322 -286 332 -285
rect 334 -281 340 -280
rect 334 -285 335 -281
rect 339 -285 340 -281
rect 334 -286 340 -285
rect 342 -281 352 -280
rect 342 -285 345 -281
rect 352 -285 353 -282
rect 357 -285 358 -282
rect 377 -281 387 -280
rect 371 -285 372 -282
rect 376 -285 377 -282
rect 384 -285 387 -281
rect 342 -286 352 -285
rect 377 -286 387 -285
rect 389 -281 395 -280
rect 389 -285 390 -281
rect 394 -285 395 -281
rect 389 -286 395 -285
rect 397 -281 407 -280
rect 397 -285 400 -281
rect 407 -285 408 -282
rect 412 -285 413 -282
rect 432 -281 442 -280
rect 426 -285 427 -282
rect 431 -285 432 -282
rect 439 -285 442 -281
rect 397 -286 407 -285
rect 432 -286 442 -285
rect 444 -281 450 -280
rect 444 -285 445 -281
rect 449 -285 450 -281
rect 444 -286 450 -285
rect 452 -281 462 -280
rect 452 -285 455 -281
rect 462 -285 463 -282
rect 467 -285 468 -282
rect 487 -281 497 -280
rect 481 -285 482 -282
rect 486 -285 487 -282
rect 494 -285 497 -281
rect 452 -286 462 -285
rect 487 -286 497 -285
rect 499 -281 505 -280
rect 499 -285 500 -281
rect 504 -285 505 -281
rect 499 -286 505 -285
rect 507 -281 517 -280
rect 507 -285 510 -281
rect 517 -285 518 -282
rect 522 -285 523 -282
rect 542 -281 552 -280
rect 536 -285 537 -282
rect 541 -285 542 -282
rect 549 -285 552 -281
rect 507 -286 517 -285
rect 542 -286 552 -285
rect 554 -281 560 -280
rect 554 -285 555 -281
rect 559 -285 560 -281
rect 554 -286 560 -285
rect 562 -281 572 -280
rect 562 -285 565 -281
rect 572 -285 573 -282
rect 577 -285 578 -282
rect 597 -281 607 -280
rect 591 -285 592 -282
rect 596 -285 597 -282
rect 604 -285 607 -281
rect 562 -286 572 -285
rect 597 -286 607 -285
rect 609 -281 615 -280
rect 609 -285 610 -281
rect 614 -285 615 -281
rect 609 -286 615 -285
rect 617 -281 627 -280
rect 617 -285 620 -281
rect 627 -285 628 -282
rect 632 -285 633 -282
rect 617 -286 627 -285
rect 212 -335 222 -334
rect 206 -338 207 -335
rect 211 -338 212 -335
rect 219 -339 222 -335
rect 212 -340 222 -339
rect 224 -335 230 -334
rect 224 -339 225 -335
rect 229 -339 230 -335
rect 224 -340 230 -339
rect 232 -335 242 -334
rect 267 -335 277 -334
rect 232 -339 235 -335
rect 242 -338 243 -335
rect 247 -338 248 -335
rect 232 -340 242 -339
rect 261 -338 262 -335
rect 266 -338 267 -335
rect 274 -339 277 -335
rect 267 -340 277 -339
rect 279 -335 285 -334
rect 279 -339 280 -335
rect 284 -339 285 -335
rect 279 -340 285 -339
rect 287 -335 297 -334
rect 322 -335 332 -334
rect 287 -339 290 -335
rect 297 -338 298 -335
rect 302 -338 303 -335
rect 287 -340 297 -339
rect 316 -338 317 -335
rect 321 -338 322 -335
rect 329 -339 332 -335
rect 322 -340 332 -339
rect 334 -335 340 -334
rect 334 -339 335 -335
rect 339 -339 340 -335
rect 334 -340 340 -339
rect 342 -335 352 -334
rect 377 -335 387 -334
rect 342 -339 345 -335
rect 352 -338 353 -335
rect 357 -338 358 -335
rect 342 -340 352 -339
rect 371 -338 372 -335
rect 376 -338 377 -335
rect 384 -339 387 -335
rect 377 -340 387 -339
rect 389 -335 395 -334
rect 389 -339 390 -335
rect 394 -339 395 -335
rect 389 -340 395 -339
rect 397 -335 407 -334
rect 432 -335 442 -334
rect 397 -339 400 -335
rect 407 -338 408 -335
rect 412 -338 413 -335
rect 397 -340 407 -339
rect 426 -338 427 -335
rect 431 -338 432 -335
rect 439 -339 442 -335
rect 432 -340 442 -339
rect 444 -335 450 -334
rect 444 -339 445 -335
rect 449 -339 450 -335
rect 444 -340 450 -339
rect 452 -335 462 -334
rect 487 -335 497 -334
rect 452 -339 455 -335
rect 462 -338 463 -335
rect 467 -338 468 -335
rect 452 -340 462 -339
rect 481 -338 482 -335
rect 486 -338 487 -335
rect 494 -339 497 -335
rect 487 -340 497 -339
rect 499 -335 505 -334
rect 499 -339 500 -335
rect 504 -339 505 -335
rect 499 -340 505 -339
rect 507 -335 517 -334
rect 542 -335 552 -334
rect 507 -339 510 -335
rect 517 -338 518 -335
rect 522 -338 523 -335
rect 507 -340 517 -339
rect 536 -338 537 -335
rect 541 -338 542 -335
rect 549 -339 552 -335
rect 542 -340 552 -339
rect 554 -335 560 -334
rect 554 -339 555 -335
rect 559 -339 560 -335
rect 554 -340 560 -339
rect 562 -335 572 -334
rect 597 -335 607 -334
rect 562 -339 565 -335
rect 572 -338 573 -335
rect 577 -338 578 -335
rect 562 -340 572 -339
rect 591 -338 592 -335
rect 596 -338 597 -335
rect 604 -339 607 -335
rect 597 -340 607 -339
rect 609 -335 615 -334
rect 609 -339 610 -335
rect 614 -339 615 -335
rect 609 -340 615 -339
rect 617 -335 627 -334
rect 617 -339 620 -335
rect 627 -338 628 -335
rect 632 -338 633 -335
rect 617 -340 627 -339
rect 212 -353 222 -352
rect 206 -357 207 -354
rect 211 -357 212 -354
rect 219 -357 222 -353
rect 212 -358 222 -357
rect 224 -353 230 -352
rect 224 -357 225 -353
rect 229 -357 230 -353
rect 224 -358 230 -357
rect 232 -353 242 -352
rect 232 -357 235 -353
rect 242 -357 243 -354
rect 247 -357 248 -354
rect 267 -353 277 -352
rect 261 -357 262 -354
rect 266 -357 267 -354
rect 274 -357 277 -353
rect 232 -358 242 -357
rect 267 -358 277 -357
rect 279 -353 285 -352
rect 279 -357 280 -353
rect 284 -357 285 -353
rect 279 -358 285 -357
rect 287 -353 297 -352
rect 287 -357 290 -353
rect 297 -357 298 -354
rect 302 -357 303 -354
rect 322 -353 332 -352
rect 316 -357 317 -354
rect 321 -357 322 -354
rect 329 -357 332 -353
rect 287 -358 297 -357
rect 322 -358 332 -357
rect 334 -353 340 -352
rect 334 -357 335 -353
rect 339 -357 340 -353
rect 334 -358 340 -357
rect 342 -353 352 -352
rect 342 -357 345 -353
rect 352 -357 353 -354
rect 357 -357 358 -354
rect 377 -353 387 -352
rect 371 -357 372 -354
rect 376 -357 377 -354
rect 384 -357 387 -353
rect 342 -358 352 -357
rect 377 -358 387 -357
rect 389 -353 395 -352
rect 389 -357 390 -353
rect 394 -357 395 -353
rect 389 -358 395 -357
rect 397 -353 407 -352
rect 397 -357 400 -353
rect 407 -357 408 -354
rect 412 -357 413 -354
rect 432 -353 442 -352
rect 426 -357 427 -354
rect 431 -357 432 -354
rect 439 -357 442 -353
rect 397 -358 407 -357
rect 432 -358 442 -357
rect 444 -353 450 -352
rect 444 -357 445 -353
rect 449 -357 450 -353
rect 444 -358 450 -357
rect 452 -353 462 -352
rect 452 -357 455 -353
rect 462 -357 463 -354
rect 467 -357 468 -354
rect 487 -353 497 -352
rect 481 -357 482 -354
rect 486 -357 487 -354
rect 494 -357 497 -353
rect 452 -358 462 -357
rect 487 -358 497 -357
rect 499 -353 505 -352
rect 499 -357 500 -353
rect 504 -357 505 -353
rect 499 -358 505 -357
rect 507 -353 517 -352
rect 507 -357 510 -353
rect 517 -357 518 -354
rect 522 -357 523 -354
rect 542 -353 552 -352
rect 536 -357 537 -354
rect 541 -357 542 -354
rect 549 -357 552 -353
rect 507 -358 517 -357
rect 542 -358 552 -357
rect 554 -353 560 -352
rect 554 -357 555 -353
rect 559 -357 560 -353
rect 554 -358 560 -357
rect 562 -353 572 -352
rect 562 -357 565 -353
rect 572 -357 573 -354
rect 577 -357 578 -354
rect 597 -353 607 -352
rect 591 -357 592 -354
rect 596 -357 597 -354
rect 604 -357 607 -353
rect 562 -358 572 -357
rect 597 -358 607 -357
rect 609 -353 615 -352
rect 609 -357 610 -353
rect 614 -357 615 -353
rect 609 -358 615 -357
rect 617 -353 627 -352
rect 617 -357 620 -353
rect 627 -357 628 -354
rect 632 -357 633 -354
rect 617 -358 627 -357
<< pdiffusion >>
rect 217 -103 218 -100
rect 224 -103 225 -100
rect 229 -103 230 -100
rect 236 -103 237 -100
rect 272 -103 273 -100
rect 279 -103 280 -100
rect 284 -103 285 -100
rect 291 -103 292 -100
rect 327 -103 328 -100
rect 334 -103 335 -100
rect 339 -103 340 -100
rect 346 -103 347 -100
rect 382 -103 383 -100
rect 389 -103 390 -100
rect 394 -103 395 -100
rect 401 -103 402 -100
rect 437 -103 438 -100
rect 444 -103 445 -100
rect 449 -103 450 -100
rect 456 -103 457 -100
rect 492 -103 493 -100
rect 499 -103 500 -100
rect 504 -103 505 -100
rect 511 -103 512 -100
rect 547 -103 548 -100
rect 554 -103 555 -100
rect 559 -103 560 -100
rect 566 -103 567 -100
rect 602 -103 603 -100
rect 609 -103 610 -100
rect 614 -103 615 -100
rect 621 -103 622 -100
rect 217 -160 218 -157
rect 224 -160 225 -157
rect 229 -160 230 -157
rect 236 -160 237 -157
rect 272 -160 273 -157
rect 279 -160 280 -157
rect 284 -160 285 -157
rect 291 -160 292 -157
rect 327 -160 328 -157
rect 334 -160 335 -157
rect 339 -160 340 -157
rect 346 -160 347 -157
rect 382 -160 383 -157
rect 389 -160 390 -157
rect 394 -160 395 -157
rect 401 -160 402 -157
rect 437 -160 438 -157
rect 444 -160 445 -157
rect 449 -160 450 -157
rect 456 -160 457 -157
rect 492 -160 493 -157
rect 499 -160 500 -157
rect 504 -160 505 -157
rect 511 -160 512 -157
rect 547 -160 548 -157
rect 554 -160 555 -157
rect 559 -160 560 -157
rect 566 -160 567 -157
rect 602 -160 603 -157
rect 609 -160 610 -157
rect 614 -160 615 -157
rect 621 -160 622 -157
rect 217 -175 218 -172
rect 224 -175 225 -172
rect 229 -175 230 -172
rect 236 -175 237 -172
rect 272 -175 273 -172
rect 279 -175 280 -172
rect 284 -175 285 -172
rect 291 -175 292 -172
rect 327 -175 328 -172
rect 334 -175 335 -172
rect 339 -175 340 -172
rect 346 -175 347 -172
rect 382 -175 383 -172
rect 389 -175 390 -172
rect 394 -175 395 -172
rect 401 -175 402 -172
rect 437 -175 438 -172
rect 444 -175 445 -172
rect 449 -175 450 -172
rect 456 -175 457 -172
rect 492 -175 493 -172
rect 499 -175 500 -172
rect 504 -175 505 -172
rect 511 -175 512 -172
rect 547 -175 548 -172
rect 554 -175 555 -172
rect 559 -175 560 -172
rect 566 -175 567 -172
rect 602 -175 603 -172
rect 609 -175 610 -172
rect 614 -175 615 -172
rect 621 -175 622 -172
rect 217 -232 218 -229
rect 224 -232 225 -229
rect 229 -232 230 -229
rect 236 -232 237 -229
rect 272 -232 273 -229
rect 279 -232 280 -229
rect 284 -232 285 -229
rect 291 -232 292 -229
rect 327 -232 328 -229
rect 334 -232 335 -229
rect 339 -232 340 -229
rect 346 -232 347 -229
rect 382 -232 383 -229
rect 389 -232 390 -229
rect 394 -232 395 -229
rect 401 -232 402 -229
rect 437 -232 438 -229
rect 444 -232 445 -229
rect 449 -232 450 -229
rect 456 -232 457 -229
rect 492 -232 493 -229
rect 499 -232 500 -229
rect 504 -232 505 -229
rect 511 -232 512 -229
rect 547 -232 548 -229
rect 554 -232 555 -229
rect 559 -232 560 -229
rect 566 -232 567 -229
rect 602 -232 603 -229
rect 609 -232 610 -229
rect 614 -232 615 -229
rect 621 -232 622 -229
rect 217 -247 218 -244
rect 224 -247 225 -244
rect 229 -247 230 -244
rect 236 -247 237 -244
rect 272 -247 273 -244
rect 279 -247 280 -244
rect 284 -247 285 -244
rect 291 -247 292 -244
rect 327 -247 328 -244
rect 334 -247 335 -244
rect 339 -247 340 -244
rect 346 -247 347 -244
rect 382 -247 383 -244
rect 389 -247 390 -244
rect 394 -247 395 -244
rect 401 -247 402 -244
rect 437 -247 438 -244
rect 444 -247 445 -244
rect 449 -247 450 -244
rect 456 -247 457 -244
rect 492 -247 493 -244
rect 499 -247 500 -244
rect 504 -247 505 -244
rect 511 -247 512 -244
rect 547 -247 548 -244
rect 554 -247 555 -244
rect 559 -247 560 -244
rect 566 -247 567 -244
rect 602 -247 603 -244
rect 609 -247 610 -244
rect 614 -247 615 -244
rect 621 -247 622 -244
rect 217 -304 218 -301
rect 224 -304 225 -301
rect 229 -304 230 -301
rect 236 -304 237 -301
rect 272 -304 273 -301
rect 279 -304 280 -301
rect 284 -304 285 -301
rect 291 -304 292 -301
rect 327 -304 328 -301
rect 334 -304 335 -301
rect 339 -304 340 -301
rect 346 -304 347 -301
rect 382 -304 383 -301
rect 389 -304 390 -301
rect 394 -304 395 -301
rect 401 -304 402 -301
rect 437 -304 438 -301
rect 444 -304 445 -301
rect 449 -304 450 -301
rect 456 -304 457 -301
rect 492 -304 493 -301
rect 499 -304 500 -301
rect 504 -304 505 -301
rect 511 -304 512 -301
rect 547 -304 548 -301
rect 554 -304 555 -301
rect 559 -304 560 -301
rect 566 -304 567 -301
rect 602 -304 603 -301
rect 609 -304 610 -301
rect 614 -304 615 -301
rect 621 -304 622 -301
rect 217 -319 218 -316
rect 224 -319 225 -316
rect 229 -319 230 -316
rect 236 -319 237 -316
rect 272 -319 273 -316
rect 279 -319 280 -316
rect 284 -319 285 -316
rect 291 -319 292 -316
rect 327 -319 328 -316
rect 334 -319 335 -316
rect 339 -319 340 -316
rect 346 -319 347 -316
rect 382 -319 383 -316
rect 389 -319 390 -316
rect 394 -319 395 -316
rect 401 -319 402 -316
rect 437 -319 438 -316
rect 444 -319 445 -316
rect 449 -319 450 -316
rect 456 -319 457 -316
rect 492 -319 493 -316
rect 499 -319 500 -316
rect 504 -319 505 -316
rect 511 -319 512 -316
rect 547 -319 548 -316
rect 554 -319 555 -316
rect 559 -319 560 -316
rect 566 -319 567 -316
rect 602 -319 603 -316
rect 609 -319 610 -316
rect 614 -319 615 -316
rect 621 -319 622 -316
rect 217 -376 218 -373
rect 224 -376 225 -373
rect 229 -376 230 -373
rect 236 -376 237 -373
rect 272 -376 273 -373
rect 279 -376 280 -373
rect 284 -376 285 -373
rect 291 -376 292 -373
rect 327 -376 328 -373
rect 334 -376 335 -373
rect 339 -376 340 -373
rect 346 -376 347 -373
rect 382 -376 383 -373
rect 389 -376 390 -373
rect 394 -376 395 -373
rect 401 -376 402 -373
rect 437 -376 438 -373
rect 444 -376 445 -373
rect 449 -376 450 -373
rect 456 -376 457 -373
rect 492 -376 493 -373
rect 499 -376 500 -373
rect 504 -376 505 -373
rect 511 -376 512 -373
rect 547 -376 548 -373
rect 554 -376 555 -373
rect 559 -376 560 -373
rect 566 -376 567 -373
rect 602 -376 603 -373
rect 609 -376 610 -373
rect 614 -376 615 -373
rect 621 -376 622 -373
<< ndcontact >>
rect 202 -123 206 -119
rect 212 -123 219 -119
rect 225 -123 229 -119
rect 235 -123 242 -119
rect 248 -123 252 -119
rect 257 -123 261 -119
rect 267 -123 274 -119
rect 280 -123 284 -119
rect 290 -123 297 -119
rect 303 -123 307 -119
rect 312 -123 316 -119
rect 322 -123 329 -119
rect 335 -123 339 -119
rect 345 -123 352 -119
rect 358 -123 362 -119
rect 367 -123 371 -119
rect 377 -123 384 -119
rect 390 -123 394 -119
rect 400 -123 407 -119
rect 413 -123 417 -119
rect 422 -123 426 -119
rect 432 -123 439 -119
rect 445 -123 449 -119
rect 455 -123 462 -119
rect 468 -123 472 -119
rect 477 -123 481 -119
rect 487 -123 494 -119
rect 500 -123 504 -119
rect 510 -123 517 -119
rect 523 -123 527 -119
rect 532 -123 536 -119
rect 542 -123 549 -119
rect 555 -123 559 -119
rect 565 -123 572 -119
rect 578 -123 582 -119
rect 587 -123 591 -119
rect 597 -123 604 -119
rect 610 -123 614 -119
rect 620 -123 627 -119
rect 633 -123 637 -119
rect 202 -141 206 -137
rect 212 -141 219 -137
rect 225 -141 229 -137
rect 235 -141 242 -137
rect 248 -141 252 -137
rect 257 -141 261 -137
rect 267 -141 274 -137
rect 280 -141 284 -137
rect 290 -141 297 -137
rect 303 -141 307 -137
rect 312 -141 316 -137
rect 322 -141 329 -137
rect 335 -141 339 -137
rect 345 -141 352 -137
rect 358 -141 362 -137
rect 367 -141 371 -137
rect 377 -141 384 -137
rect 390 -141 394 -137
rect 400 -141 407 -137
rect 413 -141 417 -137
rect 422 -141 426 -137
rect 432 -141 439 -137
rect 445 -141 449 -137
rect 455 -141 462 -137
rect 468 -141 472 -137
rect 477 -141 481 -137
rect 487 -141 494 -137
rect 500 -141 504 -137
rect 510 -141 517 -137
rect 523 -141 527 -137
rect 532 -141 536 -137
rect 542 -141 549 -137
rect 555 -141 559 -137
rect 565 -141 572 -137
rect 578 -141 582 -137
rect 587 -141 591 -137
rect 597 -141 604 -137
rect 610 -141 614 -137
rect 620 -141 627 -137
rect 633 -141 637 -137
rect 202 -195 206 -191
rect 212 -195 219 -191
rect 225 -195 229 -191
rect 235 -195 242 -191
rect 248 -195 252 -191
rect 257 -195 261 -191
rect 267 -195 274 -191
rect 280 -195 284 -191
rect 290 -195 297 -191
rect 303 -195 307 -191
rect 312 -195 316 -191
rect 322 -195 329 -191
rect 335 -195 339 -191
rect 345 -195 352 -191
rect 358 -195 362 -191
rect 367 -195 371 -191
rect 377 -195 384 -191
rect 390 -195 394 -191
rect 400 -195 407 -191
rect 413 -195 417 -191
rect 422 -195 426 -191
rect 432 -195 439 -191
rect 445 -195 449 -191
rect 455 -195 462 -191
rect 468 -195 472 -191
rect 477 -195 481 -191
rect 487 -195 494 -191
rect 500 -195 504 -191
rect 510 -195 517 -191
rect 523 -195 527 -191
rect 532 -195 536 -191
rect 542 -195 549 -191
rect 555 -195 559 -191
rect 565 -195 572 -191
rect 578 -195 582 -191
rect 587 -195 591 -191
rect 597 -195 604 -191
rect 610 -195 614 -191
rect 620 -195 627 -191
rect 633 -195 637 -191
rect 202 -213 206 -209
rect 212 -213 219 -209
rect 225 -213 229 -209
rect 235 -213 242 -209
rect 248 -213 252 -209
rect 257 -213 261 -209
rect 267 -213 274 -209
rect 280 -213 284 -209
rect 290 -213 297 -209
rect 303 -213 307 -209
rect 312 -213 316 -209
rect 322 -213 329 -209
rect 335 -213 339 -209
rect 345 -213 352 -209
rect 358 -213 362 -209
rect 367 -213 371 -209
rect 377 -213 384 -209
rect 390 -213 394 -209
rect 400 -213 407 -209
rect 413 -213 417 -209
rect 422 -213 426 -209
rect 432 -213 439 -209
rect 445 -213 449 -209
rect 455 -213 462 -209
rect 468 -213 472 -209
rect 477 -213 481 -209
rect 487 -213 494 -209
rect 500 -213 504 -209
rect 510 -213 517 -209
rect 523 -213 527 -209
rect 532 -213 536 -209
rect 542 -213 549 -209
rect 555 -213 559 -209
rect 565 -213 572 -209
rect 578 -213 582 -209
rect 587 -213 591 -209
rect 597 -213 604 -209
rect 610 -213 614 -209
rect 620 -213 627 -209
rect 633 -213 637 -209
rect 202 -267 206 -263
rect 212 -267 219 -263
rect 225 -267 229 -263
rect 235 -267 242 -263
rect 248 -267 252 -263
rect 257 -267 261 -263
rect 267 -267 274 -263
rect 280 -267 284 -263
rect 290 -267 297 -263
rect 303 -267 307 -263
rect 312 -267 316 -263
rect 322 -267 329 -263
rect 335 -267 339 -263
rect 345 -267 352 -263
rect 358 -267 362 -263
rect 367 -267 371 -263
rect 377 -267 384 -263
rect 390 -267 394 -263
rect 400 -267 407 -263
rect 413 -267 417 -263
rect 422 -267 426 -263
rect 432 -267 439 -263
rect 445 -267 449 -263
rect 455 -267 462 -263
rect 468 -267 472 -263
rect 477 -267 481 -263
rect 487 -267 494 -263
rect 500 -267 504 -263
rect 510 -267 517 -263
rect 523 -267 527 -263
rect 532 -267 536 -263
rect 542 -267 549 -263
rect 555 -267 559 -263
rect 565 -267 572 -263
rect 578 -267 582 -263
rect 587 -267 591 -263
rect 597 -267 604 -263
rect 610 -267 614 -263
rect 620 -267 627 -263
rect 633 -267 637 -263
rect 202 -285 206 -281
rect 212 -285 219 -281
rect 225 -285 229 -281
rect 235 -285 242 -281
rect 248 -285 252 -281
rect 257 -285 261 -281
rect 267 -285 274 -281
rect 280 -285 284 -281
rect 290 -285 297 -281
rect 303 -285 307 -281
rect 312 -285 316 -281
rect 322 -285 329 -281
rect 335 -285 339 -281
rect 345 -285 352 -281
rect 358 -285 362 -281
rect 367 -285 371 -281
rect 377 -285 384 -281
rect 390 -285 394 -281
rect 400 -285 407 -281
rect 413 -285 417 -281
rect 422 -285 426 -281
rect 432 -285 439 -281
rect 445 -285 449 -281
rect 455 -285 462 -281
rect 468 -285 472 -281
rect 477 -285 481 -281
rect 487 -285 494 -281
rect 500 -285 504 -281
rect 510 -285 517 -281
rect 523 -285 527 -281
rect 532 -285 536 -281
rect 542 -285 549 -281
rect 555 -285 559 -281
rect 565 -285 572 -281
rect 578 -285 582 -281
rect 587 -285 591 -281
rect 597 -285 604 -281
rect 610 -285 614 -281
rect 620 -285 627 -281
rect 633 -285 637 -281
rect 202 -339 206 -335
rect 212 -339 219 -335
rect 225 -339 229 -335
rect 235 -339 242 -335
rect 248 -339 252 -335
rect 257 -339 261 -335
rect 267 -339 274 -335
rect 280 -339 284 -335
rect 290 -339 297 -335
rect 303 -339 307 -335
rect 312 -339 316 -335
rect 322 -339 329 -335
rect 335 -339 339 -335
rect 345 -339 352 -335
rect 358 -339 362 -335
rect 367 -339 371 -335
rect 377 -339 384 -335
rect 390 -339 394 -335
rect 400 -339 407 -335
rect 413 -339 417 -335
rect 422 -339 426 -335
rect 432 -339 439 -335
rect 445 -339 449 -335
rect 455 -339 462 -335
rect 468 -339 472 -335
rect 477 -339 481 -335
rect 487 -339 494 -335
rect 500 -339 504 -335
rect 510 -339 517 -335
rect 523 -339 527 -335
rect 532 -339 536 -335
rect 542 -339 549 -335
rect 555 -339 559 -335
rect 565 -339 572 -335
rect 578 -339 582 -335
rect 587 -339 591 -335
rect 597 -339 604 -335
rect 610 -339 614 -335
rect 620 -339 627 -335
rect 633 -339 637 -335
rect 202 -357 206 -353
rect 212 -357 219 -353
rect 225 -357 229 -353
rect 235 -357 242 -353
rect 248 -357 252 -353
rect 257 -357 261 -353
rect 267 -357 274 -353
rect 280 -357 284 -353
rect 290 -357 297 -353
rect 303 -357 307 -353
rect 312 -357 316 -353
rect 322 -357 329 -353
rect 335 -357 339 -353
rect 345 -357 352 -353
rect 358 -357 362 -353
rect 367 -357 371 -353
rect 377 -357 384 -353
rect 390 -357 394 -353
rect 400 -357 407 -353
rect 413 -357 417 -353
rect 422 -357 426 -353
rect 432 -357 439 -353
rect 445 -357 449 -353
rect 455 -357 462 -353
rect 468 -357 472 -353
rect 477 -357 481 -353
rect 487 -357 494 -353
rect 500 -357 504 -353
rect 510 -357 517 -353
rect 523 -357 527 -353
rect 532 -357 536 -353
rect 542 -357 549 -353
rect 555 -357 559 -353
rect 565 -357 572 -353
rect 578 -357 582 -353
rect 587 -357 591 -353
rect 597 -357 604 -353
rect 610 -357 614 -353
rect 620 -357 627 -353
rect 633 -357 637 -353
<< pdcontact >>
rect 213 -104 217 -100
rect 225 -103 229 -99
rect 237 -104 241 -100
rect 268 -104 272 -100
rect 280 -103 284 -99
rect 292 -104 296 -100
rect 323 -104 327 -100
rect 335 -103 339 -99
rect 347 -104 351 -100
rect 378 -104 382 -100
rect 390 -103 394 -99
rect 402 -104 406 -100
rect 433 -104 437 -100
rect 445 -103 449 -99
rect 457 -104 461 -100
rect 488 -104 492 -100
rect 500 -103 504 -99
rect 512 -104 516 -100
rect 543 -104 547 -100
rect 555 -103 559 -99
rect 567 -104 571 -100
rect 598 -104 602 -100
rect 610 -103 614 -99
rect 622 -104 626 -100
rect 213 -160 217 -156
rect 225 -161 229 -157
rect 237 -160 241 -156
rect 268 -160 272 -156
rect 280 -161 284 -157
rect 292 -160 296 -156
rect 323 -160 327 -156
rect 335 -161 339 -157
rect 347 -160 351 -156
rect 378 -160 382 -156
rect 390 -161 394 -157
rect 402 -160 406 -156
rect 433 -160 437 -156
rect 445 -161 449 -157
rect 457 -160 461 -156
rect 488 -160 492 -156
rect 500 -161 504 -157
rect 512 -160 516 -156
rect 543 -160 547 -156
rect 555 -161 559 -157
rect 567 -160 571 -156
rect 598 -160 602 -156
rect 610 -161 614 -157
rect 622 -160 626 -156
rect 213 -176 217 -172
rect 225 -175 229 -171
rect 237 -176 241 -172
rect 268 -176 272 -172
rect 280 -175 284 -171
rect 292 -176 296 -172
rect 323 -176 327 -172
rect 335 -175 339 -171
rect 347 -176 351 -172
rect 378 -176 382 -172
rect 390 -175 394 -171
rect 402 -176 406 -172
rect 433 -176 437 -172
rect 445 -175 449 -171
rect 457 -176 461 -172
rect 488 -176 492 -172
rect 500 -175 504 -171
rect 512 -176 516 -172
rect 543 -176 547 -172
rect 555 -175 559 -171
rect 567 -176 571 -172
rect 598 -176 602 -172
rect 610 -175 614 -171
rect 622 -176 626 -172
rect 213 -232 217 -228
rect 225 -233 229 -229
rect 237 -232 241 -228
rect 268 -232 272 -228
rect 280 -233 284 -229
rect 292 -232 296 -228
rect 323 -232 327 -228
rect 335 -233 339 -229
rect 347 -232 351 -228
rect 378 -232 382 -228
rect 390 -233 394 -229
rect 402 -232 406 -228
rect 433 -232 437 -228
rect 445 -233 449 -229
rect 457 -232 461 -228
rect 488 -232 492 -228
rect 500 -233 504 -229
rect 512 -232 516 -228
rect 543 -232 547 -228
rect 555 -233 559 -229
rect 567 -232 571 -228
rect 598 -232 602 -228
rect 610 -233 614 -229
rect 622 -232 626 -228
rect 213 -248 217 -244
rect 225 -247 229 -243
rect 237 -248 241 -244
rect 268 -248 272 -244
rect 280 -247 284 -243
rect 292 -248 296 -244
rect 323 -248 327 -244
rect 335 -247 339 -243
rect 347 -248 351 -244
rect 378 -248 382 -244
rect 390 -247 394 -243
rect 402 -248 406 -244
rect 433 -248 437 -244
rect 445 -247 449 -243
rect 457 -248 461 -244
rect 488 -248 492 -244
rect 500 -247 504 -243
rect 512 -248 516 -244
rect 543 -248 547 -244
rect 555 -247 559 -243
rect 567 -248 571 -244
rect 598 -248 602 -244
rect 610 -247 614 -243
rect 622 -248 626 -244
rect 213 -304 217 -300
rect 225 -305 229 -301
rect 237 -304 241 -300
rect 268 -304 272 -300
rect 280 -305 284 -301
rect 292 -304 296 -300
rect 323 -304 327 -300
rect 335 -305 339 -301
rect 347 -304 351 -300
rect 378 -304 382 -300
rect 390 -305 394 -301
rect 402 -304 406 -300
rect 433 -304 437 -300
rect 445 -305 449 -301
rect 457 -304 461 -300
rect 488 -304 492 -300
rect 500 -305 504 -301
rect 512 -304 516 -300
rect 543 -304 547 -300
rect 555 -305 559 -301
rect 567 -304 571 -300
rect 598 -304 602 -300
rect 610 -305 614 -301
rect 622 -304 626 -300
rect 213 -320 217 -316
rect 225 -319 229 -315
rect 237 -320 241 -316
rect 268 -320 272 -316
rect 280 -319 284 -315
rect 292 -320 296 -316
rect 323 -320 327 -316
rect 335 -319 339 -315
rect 347 -320 351 -316
rect 378 -320 382 -316
rect 390 -319 394 -315
rect 402 -320 406 -316
rect 433 -320 437 -316
rect 445 -319 449 -315
rect 457 -320 461 -316
rect 488 -320 492 -316
rect 500 -319 504 -315
rect 512 -320 516 -316
rect 543 -320 547 -316
rect 555 -319 559 -315
rect 567 -320 571 -316
rect 598 -320 602 -316
rect 610 -319 614 -315
rect 622 -320 626 -316
rect 213 -376 217 -372
rect 225 -377 229 -373
rect 237 -376 241 -372
rect 268 -376 272 -372
rect 280 -377 284 -373
rect 292 -376 296 -372
rect 323 -376 327 -372
rect 335 -377 339 -373
rect 347 -376 351 -372
rect 378 -376 382 -372
rect 390 -377 394 -373
rect 402 -376 406 -372
rect 433 -376 437 -372
rect 445 -377 449 -373
rect 457 -376 461 -372
rect 488 -376 492 -372
rect 500 -377 504 -373
rect 512 -376 516 -372
rect 543 -376 547 -372
rect 555 -377 559 -373
rect 567 -376 571 -372
rect 598 -376 602 -372
rect 610 -377 614 -373
rect 622 -376 626 -372
<< psubstratepcontact >>
rect 215 -132 219 -128
rect 235 -132 239 -128
rect 270 -132 274 -128
rect 290 -132 294 -128
rect 325 -132 329 -128
rect 345 -132 349 -128
rect 380 -132 384 -128
rect 400 -132 404 -128
rect 435 -132 439 -128
rect 455 -132 459 -128
rect 490 -132 494 -128
rect 510 -132 514 -128
rect 545 -132 549 -128
rect 565 -132 569 -128
rect 600 -132 604 -128
rect 620 -132 624 -128
rect 215 -204 219 -200
rect 235 -204 239 -200
rect 270 -204 274 -200
rect 290 -204 294 -200
rect 325 -204 329 -200
rect 345 -204 349 -200
rect 380 -204 384 -200
rect 400 -204 404 -200
rect 435 -204 439 -200
rect 455 -204 459 -200
rect 490 -204 494 -200
rect 510 -204 514 -200
rect 545 -204 549 -200
rect 565 -204 569 -200
rect 600 -204 604 -200
rect 620 -204 624 -200
rect 215 -276 219 -272
rect 235 -276 239 -272
rect 270 -276 274 -272
rect 290 -276 294 -272
rect 325 -276 329 -272
rect 345 -276 349 -272
rect 380 -276 384 -272
rect 400 -276 404 -272
rect 435 -276 439 -272
rect 455 -276 459 -272
rect 490 -276 494 -272
rect 510 -276 514 -272
rect 545 -276 549 -272
rect 565 -276 569 -272
rect 600 -276 604 -272
rect 620 -276 624 -272
rect 215 -348 219 -344
rect 235 -348 239 -344
rect 270 -348 274 -344
rect 290 -348 294 -344
rect 325 -348 329 -344
rect 345 -348 349 -344
rect 380 -348 384 -344
rect 400 -348 404 -344
rect 435 -348 439 -344
rect 455 -348 459 -344
rect 490 -348 494 -344
rect 510 -348 514 -344
rect 545 -348 549 -344
rect 565 -348 569 -344
rect 600 -348 604 -344
rect 620 -348 624 -344
<< nsubstratencontact >>
rect 213 -96 217 -92
rect 237 -96 241 -92
rect 268 -96 272 -92
rect 292 -96 296 -92
rect 323 -96 327 -92
rect 347 -96 351 -92
rect 378 -96 382 -92
rect 402 -96 406 -92
rect 433 -96 437 -92
rect 457 -96 461 -92
rect 488 -96 492 -92
rect 512 -96 516 -92
rect 543 -96 547 -92
rect 567 -96 571 -92
rect 598 -96 602 -92
rect 622 -96 626 -92
rect 213 -168 217 -164
rect 237 -168 241 -164
rect 268 -168 272 -164
rect 292 -168 296 -164
rect 323 -168 327 -164
rect 347 -168 351 -164
rect 378 -168 382 -164
rect 402 -168 406 -164
rect 433 -168 437 -164
rect 457 -168 461 -164
rect 488 -168 492 -164
rect 512 -168 516 -164
rect 543 -168 547 -164
rect 567 -168 571 -164
rect 598 -168 602 -164
rect 622 -168 626 -164
rect 213 -240 217 -236
rect 237 -240 241 -236
rect 268 -240 272 -236
rect 292 -240 296 -236
rect 323 -240 327 -236
rect 347 -240 351 -236
rect 378 -240 382 -236
rect 402 -240 406 -236
rect 433 -240 437 -236
rect 457 -240 461 -236
rect 488 -240 492 -236
rect 512 -240 516 -236
rect 543 -240 547 -236
rect 567 -240 571 -236
rect 598 -240 602 -236
rect 622 -240 626 -236
rect 213 -312 217 -308
rect 237 -312 241 -308
rect 268 -312 272 -308
rect 292 -312 296 -308
rect 323 -312 327 -308
rect 347 -312 351 -308
rect 378 -312 382 -308
rect 402 -312 406 -308
rect 433 -312 437 -308
rect 457 -312 461 -308
rect 488 -312 492 -308
rect 512 -312 516 -308
rect 543 -312 547 -308
rect 567 -312 571 -308
rect 598 -312 602 -308
rect 622 -312 626 -308
rect 213 -384 217 -380
rect 237 -384 241 -380
rect 268 -384 272 -380
rect 292 -384 296 -380
rect 323 -384 327 -380
rect 347 -384 351 -380
rect 378 -384 382 -380
rect 402 -384 406 -380
rect 433 -384 437 -380
rect 457 -384 461 -380
rect 488 -384 492 -380
rect 512 -384 516 -380
rect 543 -384 547 -380
rect 567 -384 571 -380
rect 598 -384 602 -380
rect 622 -384 626 -380
<< polysilicon >>
rect 218 -100 224 -98
rect 230 -100 236 -98
rect 273 -100 279 -98
rect 218 -105 224 -103
rect 222 -112 224 -105
rect 207 -119 211 -114
rect 222 -118 224 -116
rect 230 -105 236 -103
rect 285 -100 291 -98
rect 328 -100 334 -98
rect 273 -105 279 -103
rect 230 -106 234 -105
rect 230 -118 232 -110
rect 207 -124 211 -122
rect 243 -119 247 -114
rect 277 -112 279 -105
rect 262 -119 266 -114
rect 277 -118 279 -116
rect 285 -105 291 -103
rect 340 -100 346 -98
rect 383 -100 389 -98
rect 328 -105 334 -103
rect 285 -106 289 -105
rect 285 -118 287 -110
rect 243 -124 247 -122
rect 262 -124 266 -122
rect 298 -119 302 -114
rect 332 -112 334 -105
rect 317 -119 321 -114
rect 332 -118 334 -116
rect 340 -105 346 -103
rect 395 -100 401 -98
rect 438 -100 444 -98
rect 383 -105 389 -103
rect 340 -106 344 -105
rect 340 -118 342 -110
rect 298 -124 302 -122
rect 317 -124 321 -122
rect 353 -119 357 -114
rect 387 -112 389 -105
rect 372 -119 376 -114
rect 387 -118 389 -116
rect 395 -105 401 -103
rect 450 -100 456 -98
rect 493 -100 499 -98
rect 438 -105 444 -103
rect 395 -106 399 -105
rect 395 -118 397 -110
rect 353 -124 357 -122
rect 372 -124 376 -122
rect 408 -119 412 -114
rect 442 -112 444 -105
rect 427 -119 431 -114
rect 442 -118 444 -116
rect 450 -105 456 -103
rect 505 -100 511 -98
rect 548 -100 554 -98
rect 493 -105 499 -103
rect 450 -106 454 -105
rect 450 -118 452 -110
rect 408 -124 412 -122
rect 427 -124 431 -122
rect 463 -119 467 -114
rect 497 -112 499 -105
rect 482 -119 486 -114
rect 497 -118 499 -116
rect 505 -105 511 -103
rect 560 -100 566 -98
rect 603 -100 609 -98
rect 548 -105 554 -103
rect 505 -106 509 -105
rect 505 -118 507 -110
rect 463 -124 467 -122
rect 482 -124 486 -122
rect 518 -119 522 -114
rect 552 -112 554 -105
rect 537 -119 541 -114
rect 552 -118 554 -116
rect 560 -105 566 -103
rect 615 -100 621 -98
rect 603 -105 609 -103
rect 560 -106 564 -105
rect 560 -118 562 -110
rect 518 -124 522 -122
rect 537 -124 541 -122
rect 573 -119 577 -114
rect 607 -112 609 -105
rect 592 -119 596 -114
rect 607 -118 609 -116
rect 615 -105 621 -103
rect 615 -106 619 -105
rect 615 -118 617 -110
rect 573 -124 577 -122
rect 592 -124 596 -122
rect 628 -119 632 -114
rect 628 -124 632 -122
rect 222 -126 224 -124
rect 230 -126 232 -124
rect 277 -126 279 -124
rect 285 -126 287 -124
rect 332 -126 334 -124
rect 340 -126 342 -124
rect 387 -126 389 -124
rect 395 -126 397 -124
rect 442 -126 444 -124
rect 450 -126 452 -124
rect 497 -126 499 -124
rect 505 -126 507 -124
rect 552 -126 554 -124
rect 560 -126 562 -124
rect 607 -126 609 -124
rect 615 -126 617 -124
rect 222 -136 224 -134
rect 230 -136 232 -134
rect 277 -136 279 -134
rect 285 -136 287 -134
rect 332 -136 334 -134
rect 340 -136 342 -134
rect 387 -136 389 -134
rect 395 -136 397 -134
rect 442 -136 444 -134
rect 450 -136 452 -134
rect 497 -136 499 -134
rect 505 -136 507 -134
rect 552 -136 554 -134
rect 560 -136 562 -134
rect 607 -136 609 -134
rect 615 -136 617 -134
rect 207 -138 211 -136
rect 207 -146 211 -141
rect 243 -138 247 -136
rect 262 -138 266 -136
rect 222 -144 224 -142
rect 222 -155 224 -148
rect 218 -157 224 -155
rect 230 -150 232 -142
rect 243 -146 247 -141
rect 262 -146 266 -141
rect 298 -138 302 -136
rect 317 -138 321 -136
rect 277 -144 279 -142
rect 230 -155 234 -154
rect 277 -155 279 -148
rect 230 -157 236 -155
rect 218 -162 224 -160
rect 273 -157 279 -155
rect 285 -150 287 -142
rect 298 -146 302 -141
rect 317 -146 321 -141
rect 353 -138 357 -136
rect 372 -138 376 -136
rect 332 -144 334 -142
rect 285 -155 289 -154
rect 332 -155 334 -148
rect 285 -157 291 -155
rect 230 -162 236 -160
rect 273 -162 279 -160
rect 328 -157 334 -155
rect 340 -150 342 -142
rect 353 -146 357 -141
rect 372 -146 376 -141
rect 408 -138 412 -136
rect 427 -138 431 -136
rect 387 -144 389 -142
rect 340 -155 344 -154
rect 387 -155 389 -148
rect 340 -157 346 -155
rect 285 -162 291 -160
rect 328 -162 334 -160
rect 383 -157 389 -155
rect 395 -150 397 -142
rect 408 -146 412 -141
rect 427 -146 431 -141
rect 463 -138 467 -136
rect 482 -138 486 -136
rect 442 -144 444 -142
rect 395 -155 399 -154
rect 442 -155 444 -148
rect 395 -157 401 -155
rect 340 -162 346 -160
rect 383 -162 389 -160
rect 438 -157 444 -155
rect 450 -150 452 -142
rect 463 -146 467 -141
rect 482 -146 486 -141
rect 518 -138 522 -136
rect 537 -138 541 -136
rect 497 -144 499 -142
rect 450 -155 454 -154
rect 497 -155 499 -148
rect 450 -157 456 -155
rect 395 -162 401 -160
rect 438 -162 444 -160
rect 493 -157 499 -155
rect 505 -150 507 -142
rect 518 -146 522 -141
rect 537 -146 541 -141
rect 573 -138 577 -136
rect 592 -138 596 -136
rect 552 -144 554 -142
rect 505 -155 509 -154
rect 552 -155 554 -148
rect 505 -157 511 -155
rect 450 -162 456 -160
rect 493 -162 499 -160
rect 548 -157 554 -155
rect 560 -150 562 -142
rect 573 -146 577 -141
rect 592 -146 596 -141
rect 628 -138 632 -136
rect 607 -144 609 -142
rect 560 -155 564 -154
rect 607 -155 609 -148
rect 560 -157 566 -155
rect 505 -162 511 -160
rect 548 -162 554 -160
rect 603 -157 609 -155
rect 615 -150 617 -142
rect 628 -146 632 -141
rect 615 -155 619 -154
rect 615 -157 621 -155
rect 560 -162 566 -160
rect 603 -162 609 -160
rect 615 -162 621 -160
rect 218 -172 224 -170
rect 230 -172 236 -170
rect 273 -172 279 -170
rect 218 -177 224 -175
rect 222 -184 224 -177
rect 207 -191 211 -186
rect 222 -190 224 -188
rect 230 -177 236 -175
rect 285 -172 291 -170
rect 328 -172 334 -170
rect 273 -177 279 -175
rect 230 -178 234 -177
rect 230 -190 232 -182
rect 207 -196 211 -194
rect 243 -191 247 -186
rect 277 -184 279 -177
rect 262 -191 266 -186
rect 277 -190 279 -188
rect 285 -177 291 -175
rect 340 -172 346 -170
rect 383 -172 389 -170
rect 328 -177 334 -175
rect 285 -178 289 -177
rect 285 -190 287 -182
rect 243 -196 247 -194
rect 262 -196 266 -194
rect 298 -191 302 -186
rect 332 -184 334 -177
rect 317 -191 321 -186
rect 332 -190 334 -188
rect 340 -177 346 -175
rect 395 -172 401 -170
rect 438 -172 444 -170
rect 383 -177 389 -175
rect 340 -178 344 -177
rect 340 -190 342 -182
rect 298 -196 302 -194
rect 317 -196 321 -194
rect 353 -191 357 -186
rect 387 -184 389 -177
rect 372 -191 376 -186
rect 387 -190 389 -188
rect 395 -177 401 -175
rect 450 -172 456 -170
rect 493 -172 499 -170
rect 438 -177 444 -175
rect 395 -178 399 -177
rect 395 -190 397 -182
rect 353 -196 357 -194
rect 372 -196 376 -194
rect 408 -191 412 -186
rect 442 -184 444 -177
rect 427 -191 431 -186
rect 442 -190 444 -188
rect 450 -177 456 -175
rect 505 -172 511 -170
rect 548 -172 554 -170
rect 493 -177 499 -175
rect 450 -178 454 -177
rect 450 -190 452 -182
rect 408 -196 412 -194
rect 427 -196 431 -194
rect 463 -191 467 -186
rect 497 -184 499 -177
rect 482 -191 486 -186
rect 497 -190 499 -188
rect 505 -177 511 -175
rect 560 -172 566 -170
rect 603 -172 609 -170
rect 548 -177 554 -175
rect 505 -178 509 -177
rect 505 -190 507 -182
rect 463 -196 467 -194
rect 482 -196 486 -194
rect 518 -191 522 -186
rect 552 -184 554 -177
rect 537 -191 541 -186
rect 552 -190 554 -188
rect 560 -177 566 -175
rect 615 -172 621 -170
rect 603 -177 609 -175
rect 560 -178 564 -177
rect 560 -190 562 -182
rect 518 -196 522 -194
rect 537 -196 541 -194
rect 573 -191 577 -186
rect 607 -184 609 -177
rect 592 -191 596 -186
rect 607 -190 609 -188
rect 615 -177 621 -175
rect 615 -178 619 -177
rect 615 -190 617 -182
rect 573 -196 577 -194
rect 592 -196 596 -194
rect 628 -191 632 -186
rect 628 -196 632 -194
rect 222 -198 224 -196
rect 230 -198 232 -196
rect 277 -198 279 -196
rect 285 -198 287 -196
rect 332 -198 334 -196
rect 340 -198 342 -196
rect 387 -198 389 -196
rect 395 -198 397 -196
rect 442 -198 444 -196
rect 450 -198 452 -196
rect 497 -198 499 -196
rect 505 -198 507 -196
rect 552 -198 554 -196
rect 560 -198 562 -196
rect 607 -198 609 -196
rect 615 -198 617 -196
rect 222 -208 224 -206
rect 230 -208 232 -206
rect 277 -208 279 -206
rect 285 -208 287 -206
rect 332 -208 334 -206
rect 340 -208 342 -206
rect 387 -208 389 -206
rect 395 -208 397 -206
rect 442 -208 444 -206
rect 450 -208 452 -206
rect 497 -208 499 -206
rect 505 -208 507 -206
rect 552 -208 554 -206
rect 560 -208 562 -206
rect 607 -208 609 -206
rect 615 -208 617 -206
rect 207 -210 211 -208
rect 207 -218 211 -213
rect 243 -210 247 -208
rect 262 -210 266 -208
rect 222 -216 224 -214
rect 222 -227 224 -220
rect 218 -229 224 -227
rect 230 -222 232 -214
rect 243 -218 247 -213
rect 262 -218 266 -213
rect 298 -210 302 -208
rect 317 -210 321 -208
rect 277 -216 279 -214
rect 230 -227 234 -226
rect 277 -227 279 -220
rect 230 -229 236 -227
rect 218 -234 224 -232
rect 273 -229 279 -227
rect 285 -222 287 -214
rect 298 -218 302 -213
rect 317 -218 321 -213
rect 353 -210 357 -208
rect 372 -210 376 -208
rect 332 -216 334 -214
rect 285 -227 289 -226
rect 332 -227 334 -220
rect 285 -229 291 -227
rect 230 -234 236 -232
rect 273 -234 279 -232
rect 328 -229 334 -227
rect 340 -222 342 -214
rect 353 -218 357 -213
rect 372 -218 376 -213
rect 408 -210 412 -208
rect 427 -210 431 -208
rect 387 -216 389 -214
rect 340 -227 344 -226
rect 387 -227 389 -220
rect 340 -229 346 -227
rect 285 -234 291 -232
rect 328 -234 334 -232
rect 383 -229 389 -227
rect 395 -222 397 -214
rect 408 -218 412 -213
rect 427 -218 431 -213
rect 463 -210 467 -208
rect 482 -210 486 -208
rect 442 -216 444 -214
rect 395 -227 399 -226
rect 442 -227 444 -220
rect 395 -229 401 -227
rect 340 -234 346 -232
rect 383 -234 389 -232
rect 438 -229 444 -227
rect 450 -222 452 -214
rect 463 -218 467 -213
rect 482 -218 486 -213
rect 518 -210 522 -208
rect 537 -210 541 -208
rect 497 -216 499 -214
rect 450 -227 454 -226
rect 497 -227 499 -220
rect 450 -229 456 -227
rect 395 -234 401 -232
rect 438 -234 444 -232
rect 493 -229 499 -227
rect 505 -222 507 -214
rect 518 -218 522 -213
rect 537 -218 541 -213
rect 573 -210 577 -208
rect 592 -210 596 -208
rect 552 -216 554 -214
rect 505 -227 509 -226
rect 552 -227 554 -220
rect 505 -229 511 -227
rect 450 -234 456 -232
rect 493 -234 499 -232
rect 548 -229 554 -227
rect 560 -222 562 -214
rect 573 -218 577 -213
rect 592 -218 596 -213
rect 628 -210 632 -208
rect 607 -216 609 -214
rect 560 -227 564 -226
rect 607 -227 609 -220
rect 560 -229 566 -227
rect 505 -234 511 -232
rect 548 -234 554 -232
rect 603 -229 609 -227
rect 615 -222 617 -214
rect 628 -218 632 -213
rect 615 -227 619 -226
rect 615 -229 621 -227
rect 560 -234 566 -232
rect 603 -234 609 -232
rect 615 -234 621 -232
rect 218 -244 224 -242
rect 230 -244 236 -242
rect 273 -244 279 -242
rect 218 -249 224 -247
rect 222 -256 224 -249
rect 207 -263 211 -258
rect 222 -262 224 -260
rect 230 -249 236 -247
rect 285 -244 291 -242
rect 328 -244 334 -242
rect 273 -249 279 -247
rect 230 -250 234 -249
rect 230 -262 232 -254
rect 207 -268 211 -266
rect 243 -263 247 -258
rect 277 -256 279 -249
rect 262 -263 266 -258
rect 277 -262 279 -260
rect 285 -249 291 -247
rect 340 -244 346 -242
rect 383 -244 389 -242
rect 328 -249 334 -247
rect 285 -250 289 -249
rect 285 -262 287 -254
rect 243 -268 247 -266
rect 262 -268 266 -266
rect 298 -263 302 -258
rect 332 -256 334 -249
rect 317 -263 321 -258
rect 332 -262 334 -260
rect 340 -249 346 -247
rect 395 -244 401 -242
rect 438 -244 444 -242
rect 383 -249 389 -247
rect 340 -250 344 -249
rect 340 -262 342 -254
rect 298 -268 302 -266
rect 317 -268 321 -266
rect 353 -263 357 -258
rect 387 -256 389 -249
rect 372 -263 376 -258
rect 387 -262 389 -260
rect 395 -249 401 -247
rect 450 -244 456 -242
rect 493 -244 499 -242
rect 438 -249 444 -247
rect 395 -250 399 -249
rect 395 -262 397 -254
rect 353 -268 357 -266
rect 372 -268 376 -266
rect 408 -263 412 -258
rect 442 -256 444 -249
rect 427 -263 431 -258
rect 442 -262 444 -260
rect 450 -249 456 -247
rect 505 -244 511 -242
rect 548 -244 554 -242
rect 493 -249 499 -247
rect 450 -250 454 -249
rect 450 -262 452 -254
rect 408 -268 412 -266
rect 427 -268 431 -266
rect 463 -263 467 -258
rect 497 -256 499 -249
rect 482 -263 486 -258
rect 497 -262 499 -260
rect 505 -249 511 -247
rect 560 -244 566 -242
rect 603 -244 609 -242
rect 548 -249 554 -247
rect 505 -250 509 -249
rect 505 -262 507 -254
rect 463 -268 467 -266
rect 482 -268 486 -266
rect 518 -263 522 -258
rect 552 -256 554 -249
rect 537 -263 541 -258
rect 552 -262 554 -260
rect 560 -249 566 -247
rect 615 -244 621 -242
rect 603 -249 609 -247
rect 560 -250 564 -249
rect 560 -262 562 -254
rect 518 -268 522 -266
rect 537 -268 541 -266
rect 573 -263 577 -258
rect 607 -256 609 -249
rect 592 -263 596 -258
rect 607 -262 609 -260
rect 615 -249 621 -247
rect 615 -250 619 -249
rect 615 -262 617 -254
rect 573 -268 577 -266
rect 592 -268 596 -266
rect 628 -263 632 -258
rect 628 -268 632 -266
rect 222 -270 224 -268
rect 230 -270 232 -268
rect 277 -270 279 -268
rect 285 -270 287 -268
rect 332 -270 334 -268
rect 340 -270 342 -268
rect 387 -270 389 -268
rect 395 -270 397 -268
rect 442 -270 444 -268
rect 450 -270 452 -268
rect 497 -270 499 -268
rect 505 -270 507 -268
rect 552 -270 554 -268
rect 560 -270 562 -268
rect 607 -270 609 -268
rect 615 -270 617 -268
rect 222 -280 224 -278
rect 230 -280 232 -278
rect 277 -280 279 -278
rect 285 -280 287 -278
rect 332 -280 334 -278
rect 340 -280 342 -278
rect 387 -280 389 -278
rect 395 -280 397 -278
rect 442 -280 444 -278
rect 450 -280 452 -278
rect 497 -280 499 -278
rect 505 -280 507 -278
rect 552 -280 554 -278
rect 560 -280 562 -278
rect 607 -280 609 -278
rect 615 -280 617 -278
rect 207 -282 211 -280
rect 207 -290 211 -285
rect 243 -282 247 -280
rect 262 -282 266 -280
rect 222 -288 224 -286
rect 222 -299 224 -292
rect 218 -301 224 -299
rect 230 -294 232 -286
rect 243 -290 247 -285
rect 262 -290 266 -285
rect 298 -282 302 -280
rect 317 -282 321 -280
rect 277 -288 279 -286
rect 230 -299 234 -298
rect 277 -299 279 -292
rect 230 -301 236 -299
rect 218 -306 224 -304
rect 273 -301 279 -299
rect 285 -294 287 -286
rect 298 -290 302 -285
rect 317 -290 321 -285
rect 353 -282 357 -280
rect 372 -282 376 -280
rect 332 -288 334 -286
rect 285 -299 289 -298
rect 332 -299 334 -292
rect 285 -301 291 -299
rect 230 -306 236 -304
rect 273 -306 279 -304
rect 328 -301 334 -299
rect 340 -294 342 -286
rect 353 -290 357 -285
rect 372 -290 376 -285
rect 408 -282 412 -280
rect 427 -282 431 -280
rect 387 -288 389 -286
rect 340 -299 344 -298
rect 387 -299 389 -292
rect 340 -301 346 -299
rect 285 -306 291 -304
rect 328 -306 334 -304
rect 383 -301 389 -299
rect 395 -294 397 -286
rect 408 -290 412 -285
rect 427 -290 431 -285
rect 463 -282 467 -280
rect 482 -282 486 -280
rect 442 -288 444 -286
rect 395 -299 399 -298
rect 442 -299 444 -292
rect 395 -301 401 -299
rect 340 -306 346 -304
rect 383 -306 389 -304
rect 438 -301 444 -299
rect 450 -294 452 -286
rect 463 -290 467 -285
rect 482 -290 486 -285
rect 518 -282 522 -280
rect 537 -282 541 -280
rect 497 -288 499 -286
rect 450 -299 454 -298
rect 497 -299 499 -292
rect 450 -301 456 -299
rect 395 -306 401 -304
rect 438 -306 444 -304
rect 493 -301 499 -299
rect 505 -294 507 -286
rect 518 -290 522 -285
rect 537 -290 541 -285
rect 573 -282 577 -280
rect 592 -282 596 -280
rect 552 -288 554 -286
rect 505 -299 509 -298
rect 552 -299 554 -292
rect 505 -301 511 -299
rect 450 -306 456 -304
rect 493 -306 499 -304
rect 548 -301 554 -299
rect 560 -294 562 -286
rect 573 -290 577 -285
rect 592 -290 596 -285
rect 628 -282 632 -280
rect 607 -288 609 -286
rect 560 -299 564 -298
rect 607 -299 609 -292
rect 560 -301 566 -299
rect 505 -306 511 -304
rect 548 -306 554 -304
rect 603 -301 609 -299
rect 615 -294 617 -286
rect 628 -290 632 -285
rect 615 -299 619 -298
rect 615 -301 621 -299
rect 560 -306 566 -304
rect 603 -306 609 -304
rect 615 -306 621 -304
rect 218 -316 224 -314
rect 230 -316 236 -314
rect 273 -316 279 -314
rect 218 -321 224 -319
rect 222 -328 224 -321
rect 207 -335 211 -330
rect 222 -334 224 -332
rect 230 -321 236 -319
rect 285 -316 291 -314
rect 328 -316 334 -314
rect 273 -321 279 -319
rect 230 -322 234 -321
rect 230 -334 232 -326
rect 207 -340 211 -338
rect 243 -335 247 -330
rect 277 -328 279 -321
rect 262 -335 266 -330
rect 277 -334 279 -332
rect 285 -321 291 -319
rect 340 -316 346 -314
rect 383 -316 389 -314
rect 328 -321 334 -319
rect 285 -322 289 -321
rect 285 -334 287 -326
rect 243 -340 247 -338
rect 262 -340 266 -338
rect 298 -335 302 -330
rect 332 -328 334 -321
rect 317 -335 321 -330
rect 332 -334 334 -332
rect 340 -321 346 -319
rect 395 -316 401 -314
rect 438 -316 444 -314
rect 383 -321 389 -319
rect 340 -322 344 -321
rect 340 -334 342 -326
rect 298 -340 302 -338
rect 317 -340 321 -338
rect 353 -335 357 -330
rect 387 -328 389 -321
rect 372 -335 376 -330
rect 387 -334 389 -332
rect 395 -321 401 -319
rect 450 -316 456 -314
rect 493 -316 499 -314
rect 438 -321 444 -319
rect 395 -322 399 -321
rect 395 -334 397 -326
rect 353 -340 357 -338
rect 372 -340 376 -338
rect 408 -335 412 -330
rect 442 -328 444 -321
rect 427 -335 431 -330
rect 442 -334 444 -332
rect 450 -321 456 -319
rect 505 -316 511 -314
rect 548 -316 554 -314
rect 493 -321 499 -319
rect 450 -322 454 -321
rect 450 -334 452 -326
rect 408 -340 412 -338
rect 427 -340 431 -338
rect 463 -335 467 -330
rect 497 -328 499 -321
rect 482 -335 486 -330
rect 497 -334 499 -332
rect 505 -321 511 -319
rect 560 -316 566 -314
rect 603 -316 609 -314
rect 548 -321 554 -319
rect 505 -322 509 -321
rect 505 -334 507 -326
rect 463 -340 467 -338
rect 482 -340 486 -338
rect 518 -335 522 -330
rect 552 -328 554 -321
rect 537 -335 541 -330
rect 552 -334 554 -332
rect 560 -321 566 -319
rect 615 -316 621 -314
rect 603 -321 609 -319
rect 560 -322 564 -321
rect 560 -334 562 -326
rect 518 -340 522 -338
rect 537 -340 541 -338
rect 573 -335 577 -330
rect 607 -328 609 -321
rect 592 -335 596 -330
rect 607 -334 609 -332
rect 615 -321 621 -319
rect 615 -322 619 -321
rect 615 -334 617 -326
rect 573 -340 577 -338
rect 592 -340 596 -338
rect 628 -335 632 -330
rect 628 -340 632 -338
rect 222 -342 224 -340
rect 230 -342 232 -340
rect 277 -342 279 -340
rect 285 -342 287 -340
rect 332 -342 334 -340
rect 340 -342 342 -340
rect 387 -342 389 -340
rect 395 -342 397 -340
rect 442 -342 444 -340
rect 450 -342 452 -340
rect 497 -342 499 -340
rect 505 -342 507 -340
rect 552 -342 554 -340
rect 560 -342 562 -340
rect 607 -342 609 -340
rect 615 -342 617 -340
rect 222 -352 224 -350
rect 230 -352 232 -350
rect 277 -352 279 -350
rect 285 -352 287 -350
rect 332 -352 334 -350
rect 340 -352 342 -350
rect 387 -352 389 -350
rect 395 -352 397 -350
rect 442 -352 444 -350
rect 450 -352 452 -350
rect 497 -352 499 -350
rect 505 -352 507 -350
rect 552 -352 554 -350
rect 560 -352 562 -350
rect 607 -352 609 -350
rect 615 -352 617 -350
rect 207 -354 211 -352
rect 207 -362 211 -357
rect 243 -354 247 -352
rect 262 -354 266 -352
rect 222 -360 224 -358
rect 222 -371 224 -364
rect 218 -373 224 -371
rect 230 -366 232 -358
rect 243 -362 247 -357
rect 262 -362 266 -357
rect 298 -354 302 -352
rect 317 -354 321 -352
rect 277 -360 279 -358
rect 230 -371 234 -370
rect 277 -371 279 -364
rect 230 -373 236 -371
rect 218 -378 224 -376
rect 273 -373 279 -371
rect 285 -366 287 -358
rect 298 -362 302 -357
rect 317 -362 321 -357
rect 353 -354 357 -352
rect 372 -354 376 -352
rect 332 -360 334 -358
rect 285 -371 289 -370
rect 332 -371 334 -364
rect 285 -373 291 -371
rect 230 -378 236 -376
rect 273 -378 279 -376
rect 328 -373 334 -371
rect 340 -366 342 -358
rect 353 -362 357 -357
rect 372 -362 376 -357
rect 408 -354 412 -352
rect 427 -354 431 -352
rect 387 -360 389 -358
rect 340 -371 344 -370
rect 387 -371 389 -364
rect 340 -373 346 -371
rect 285 -378 291 -376
rect 328 -378 334 -376
rect 383 -373 389 -371
rect 395 -366 397 -358
rect 408 -362 412 -357
rect 427 -362 431 -357
rect 463 -354 467 -352
rect 482 -354 486 -352
rect 442 -360 444 -358
rect 395 -371 399 -370
rect 442 -371 444 -364
rect 395 -373 401 -371
rect 340 -378 346 -376
rect 383 -378 389 -376
rect 438 -373 444 -371
rect 450 -366 452 -358
rect 463 -362 467 -357
rect 482 -362 486 -357
rect 518 -354 522 -352
rect 537 -354 541 -352
rect 497 -360 499 -358
rect 450 -371 454 -370
rect 497 -371 499 -364
rect 450 -373 456 -371
rect 395 -378 401 -376
rect 438 -378 444 -376
rect 493 -373 499 -371
rect 505 -366 507 -358
rect 518 -362 522 -357
rect 537 -362 541 -357
rect 573 -354 577 -352
rect 592 -354 596 -352
rect 552 -360 554 -358
rect 505 -371 509 -370
rect 552 -371 554 -364
rect 505 -373 511 -371
rect 450 -378 456 -376
rect 493 -378 499 -376
rect 548 -373 554 -371
rect 560 -366 562 -358
rect 573 -362 577 -357
rect 592 -362 596 -357
rect 628 -354 632 -352
rect 607 -360 609 -358
rect 560 -371 564 -370
rect 607 -371 609 -364
rect 560 -373 566 -371
rect 505 -378 511 -376
rect 548 -378 554 -376
rect 603 -373 609 -371
rect 615 -366 617 -358
rect 628 -362 632 -357
rect 615 -371 619 -370
rect 615 -373 621 -371
rect 560 -378 566 -376
rect 603 -378 609 -376
rect 615 -378 621 -376
<< polycontact >>
rect 207 -114 211 -110
rect 220 -116 224 -112
rect 230 -110 234 -106
rect 243 -114 247 -110
rect 262 -114 266 -110
rect 275 -116 279 -112
rect 285 -110 289 -106
rect 298 -114 302 -110
rect 317 -114 321 -110
rect 330 -116 334 -112
rect 340 -110 344 -106
rect 353 -114 357 -110
rect 372 -114 376 -110
rect 385 -116 389 -112
rect 395 -110 399 -106
rect 408 -114 412 -110
rect 427 -114 431 -110
rect 440 -116 444 -112
rect 450 -110 454 -106
rect 463 -114 467 -110
rect 482 -114 486 -110
rect 495 -116 499 -112
rect 505 -110 509 -106
rect 518 -114 522 -110
rect 537 -114 541 -110
rect 550 -116 554 -112
rect 560 -110 564 -106
rect 573 -114 577 -110
rect 592 -114 596 -110
rect 605 -116 609 -112
rect 615 -110 619 -106
rect 628 -114 632 -110
rect 207 -150 211 -146
rect 220 -148 224 -144
rect 243 -150 247 -146
rect 262 -150 266 -146
rect 275 -148 279 -144
rect 230 -154 234 -150
rect 298 -150 302 -146
rect 317 -150 321 -146
rect 330 -148 334 -144
rect 285 -154 289 -150
rect 353 -150 357 -146
rect 372 -150 376 -146
rect 385 -148 389 -144
rect 340 -154 344 -150
rect 408 -150 412 -146
rect 427 -150 431 -146
rect 440 -148 444 -144
rect 395 -154 399 -150
rect 463 -150 467 -146
rect 482 -150 486 -146
rect 495 -148 499 -144
rect 450 -154 454 -150
rect 518 -150 522 -146
rect 537 -150 541 -146
rect 550 -148 554 -144
rect 505 -154 509 -150
rect 573 -150 577 -146
rect 592 -150 596 -146
rect 605 -148 609 -144
rect 560 -154 564 -150
rect 628 -150 632 -146
rect 615 -154 619 -150
rect 207 -186 211 -182
rect 220 -188 224 -184
rect 230 -182 234 -178
rect 243 -186 247 -182
rect 262 -186 266 -182
rect 275 -188 279 -184
rect 285 -182 289 -178
rect 298 -186 302 -182
rect 317 -186 321 -182
rect 330 -188 334 -184
rect 340 -182 344 -178
rect 353 -186 357 -182
rect 372 -186 376 -182
rect 385 -188 389 -184
rect 395 -182 399 -178
rect 408 -186 412 -182
rect 427 -186 431 -182
rect 440 -188 444 -184
rect 450 -182 454 -178
rect 463 -186 467 -182
rect 482 -186 486 -182
rect 495 -188 499 -184
rect 505 -182 509 -178
rect 518 -186 522 -182
rect 537 -186 541 -182
rect 550 -188 554 -184
rect 560 -182 564 -178
rect 573 -186 577 -182
rect 592 -186 596 -182
rect 605 -188 609 -184
rect 615 -182 619 -178
rect 628 -186 632 -182
rect 207 -222 211 -218
rect 220 -220 224 -216
rect 243 -222 247 -218
rect 262 -222 266 -218
rect 275 -220 279 -216
rect 230 -226 234 -222
rect 298 -222 302 -218
rect 317 -222 321 -218
rect 330 -220 334 -216
rect 285 -226 289 -222
rect 353 -222 357 -218
rect 372 -222 376 -218
rect 385 -220 389 -216
rect 340 -226 344 -222
rect 408 -222 412 -218
rect 427 -222 431 -218
rect 440 -220 444 -216
rect 395 -226 399 -222
rect 463 -222 467 -218
rect 482 -222 486 -218
rect 495 -220 499 -216
rect 450 -226 454 -222
rect 518 -222 522 -218
rect 537 -222 541 -218
rect 550 -220 554 -216
rect 505 -226 509 -222
rect 573 -222 577 -218
rect 592 -222 596 -218
rect 605 -220 609 -216
rect 560 -226 564 -222
rect 628 -222 632 -218
rect 615 -226 619 -222
rect 207 -258 211 -254
rect 220 -260 224 -256
rect 230 -254 234 -250
rect 243 -258 247 -254
rect 262 -258 266 -254
rect 275 -260 279 -256
rect 285 -254 289 -250
rect 298 -258 302 -254
rect 317 -258 321 -254
rect 330 -260 334 -256
rect 340 -254 344 -250
rect 353 -258 357 -254
rect 372 -258 376 -254
rect 385 -260 389 -256
rect 395 -254 399 -250
rect 408 -258 412 -254
rect 427 -258 431 -254
rect 440 -260 444 -256
rect 450 -254 454 -250
rect 463 -258 467 -254
rect 482 -258 486 -254
rect 495 -260 499 -256
rect 505 -254 509 -250
rect 518 -258 522 -254
rect 537 -258 541 -254
rect 550 -260 554 -256
rect 560 -254 564 -250
rect 573 -258 577 -254
rect 592 -258 596 -254
rect 605 -260 609 -256
rect 615 -254 619 -250
rect 628 -258 632 -254
rect 207 -294 211 -290
rect 220 -292 224 -288
rect 243 -294 247 -290
rect 262 -294 266 -290
rect 275 -292 279 -288
rect 230 -298 234 -294
rect 298 -294 302 -290
rect 317 -294 321 -290
rect 330 -292 334 -288
rect 285 -298 289 -294
rect 353 -294 357 -290
rect 372 -294 376 -290
rect 385 -292 389 -288
rect 340 -298 344 -294
rect 408 -294 412 -290
rect 427 -294 431 -290
rect 440 -292 444 -288
rect 395 -298 399 -294
rect 463 -294 467 -290
rect 482 -294 486 -290
rect 495 -292 499 -288
rect 450 -298 454 -294
rect 518 -294 522 -290
rect 537 -294 541 -290
rect 550 -292 554 -288
rect 505 -298 509 -294
rect 573 -294 577 -290
rect 592 -294 596 -290
rect 605 -292 609 -288
rect 560 -298 564 -294
rect 628 -294 632 -290
rect 615 -298 619 -294
rect 207 -330 211 -326
rect 220 -332 224 -328
rect 230 -326 234 -322
rect 243 -330 247 -326
rect 262 -330 266 -326
rect 275 -332 279 -328
rect 285 -326 289 -322
rect 298 -330 302 -326
rect 317 -330 321 -326
rect 330 -332 334 -328
rect 340 -326 344 -322
rect 353 -330 357 -326
rect 372 -330 376 -326
rect 385 -332 389 -328
rect 395 -326 399 -322
rect 408 -330 412 -326
rect 427 -330 431 -326
rect 440 -332 444 -328
rect 450 -326 454 -322
rect 463 -330 467 -326
rect 482 -330 486 -326
rect 495 -332 499 -328
rect 505 -326 509 -322
rect 518 -330 522 -326
rect 537 -330 541 -326
rect 550 -332 554 -328
rect 560 -326 564 -322
rect 573 -330 577 -326
rect 592 -330 596 -326
rect 605 -332 609 -328
rect 615 -326 619 -322
rect 628 -330 632 -326
rect 207 -366 211 -362
rect 220 -364 224 -360
rect 243 -366 247 -362
rect 262 -366 266 -362
rect 275 -364 279 -360
rect 230 -370 234 -366
rect 298 -366 302 -362
rect 317 -366 321 -362
rect 330 -364 334 -360
rect 285 -370 289 -366
rect 353 -366 357 -362
rect 372 -366 376 -362
rect 385 -364 389 -360
rect 340 -370 344 -366
rect 408 -366 412 -362
rect 427 -366 431 -362
rect 440 -364 444 -360
rect 395 -370 399 -366
rect 463 -366 467 -362
rect 482 -366 486 -362
rect 495 -364 499 -360
rect 450 -370 454 -366
rect 518 -366 522 -362
rect 537 -366 541 -362
rect 550 -364 554 -360
rect 505 -370 509 -366
rect 573 -366 577 -362
rect 592 -366 596 -362
rect 605 -364 609 -360
rect 560 -370 564 -366
rect 628 -366 632 -362
rect 615 -370 619 -366
<< metal1 >>
rect 201 -119 204 -92
rect 217 -96 225 -92
rect 229 -96 237 -92
rect 225 -99 229 -96
rect 214 -106 217 -104
rect 214 -109 230 -106
rect 214 -119 217 -109
rect 237 -113 240 -104
rect 224 -116 240 -113
rect 237 -119 240 -116
rect 250 -119 253 -92
rect 201 -123 202 -119
rect 252 -123 253 -119
rect 201 -137 204 -123
rect 225 -128 229 -123
rect 219 -132 225 -128
rect 229 -132 235 -128
rect 225 -137 229 -132
rect 250 -137 253 -123
rect 201 -141 202 -137
rect 252 -141 253 -137
rect 201 -191 204 -141
rect 214 -151 217 -141
rect 237 -144 240 -141
rect 224 -147 240 -144
rect 214 -154 230 -151
rect 214 -156 217 -154
rect 237 -156 240 -147
rect 225 -164 229 -161
rect 217 -168 225 -164
rect 229 -168 237 -164
rect 225 -171 229 -168
rect 214 -178 217 -176
rect 214 -181 230 -178
rect 214 -191 217 -181
rect 237 -185 240 -176
rect 224 -188 240 -185
rect 237 -191 240 -188
rect 250 -191 253 -141
rect 201 -195 202 -191
rect 252 -195 253 -191
rect 201 -209 204 -195
rect 225 -200 229 -195
rect 219 -204 225 -200
rect 229 -204 235 -200
rect 225 -209 229 -204
rect 250 -209 253 -195
rect 201 -213 202 -209
rect 252 -213 253 -209
rect 201 -263 204 -213
rect 214 -223 217 -213
rect 237 -216 240 -213
rect 224 -219 240 -216
rect 214 -226 230 -223
rect 214 -228 217 -226
rect 237 -228 240 -219
rect 225 -236 229 -233
rect 217 -240 225 -236
rect 229 -240 237 -236
rect 225 -243 229 -240
rect 214 -250 217 -248
rect 214 -253 230 -250
rect 214 -263 217 -253
rect 237 -257 240 -248
rect 224 -260 240 -257
rect 237 -263 240 -260
rect 250 -263 253 -213
rect 201 -267 202 -263
rect 252 -267 253 -263
rect 201 -281 204 -267
rect 225 -272 229 -267
rect 219 -276 225 -272
rect 229 -276 235 -272
rect 225 -281 229 -276
rect 250 -281 253 -267
rect 201 -285 202 -281
rect 252 -285 253 -281
rect 201 -335 204 -285
rect 214 -295 217 -285
rect 237 -288 240 -285
rect 224 -291 240 -288
rect 214 -298 230 -295
rect 214 -300 217 -298
rect 237 -300 240 -291
rect 225 -308 229 -305
rect 217 -312 225 -308
rect 229 -312 237 -308
rect 225 -315 229 -312
rect 214 -322 217 -320
rect 214 -325 230 -322
rect 214 -335 217 -325
rect 237 -329 240 -320
rect 224 -332 240 -329
rect 237 -335 240 -332
rect 250 -335 253 -285
rect 201 -339 202 -335
rect 252 -339 253 -335
rect 201 -353 204 -339
rect 225 -344 229 -339
rect 219 -348 225 -344
rect 229 -348 235 -344
rect 225 -353 229 -348
rect 250 -353 253 -339
rect 201 -357 202 -353
rect 252 -357 253 -353
rect 201 -387 204 -357
rect 214 -367 217 -357
rect 237 -360 240 -357
rect 224 -363 240 -360
rect 214 -370 230 -367
rect 214 -372 217 -370
rect 237 -372 240 -363
rect 225 -380 229 -377
rect 217 -384 225 -380
rect 229 -384 237 -380
rect 225 -387 229 -384
rect 250 -387 253 -357
rect 256 -119 259 -92
rect 272 -96 280 -92
rect 284 -96 292 -92
rect 280 -99 284 -96
rect 269 -106 272 -104
rect 269 -109 285 -106
rect 269 -119 272 -109
rect 292 -113 295 -104
rect 279 -116 295 -113
rect 292 -119 295 -116
rect 305 -119 308 -92
rect 256 -123 257 -119
rect 307 -123 308 -119
rect 256 -137 259 -123
rect 280 -128 284 -123
rect 274 -132 280 -128
rect 284 -132 290 -128
rect 280 -137 284 -132
rect 305 -137 308 -123
rect 256 -141 257 -137
rect 307 -141 308 -137
rect 256 -191 259 -141
rect 269 -151 272 -141
rect 292 -144 295 -141
rect 279 -147 295 -144
rect 269 -154 285 -151
rect 269 -156 272 -154
rect 292 -156 295 -147
rect 280 -164 284 -161
rect 272 -168 280 -164
rect 284 -168 292 -164
rect 280 -171 284 -168
rect 269 -178 272 -176
rect 269 -181 285 -178
rect 269 -191 272 -181
rect 292 -185 295 -176
rect 279 -188 295 -185
rect 292 -191 295 -188
rect 305 -191 308 -141
rect 256 -195 257 -191
rect 307 -195 308 -191
rect 256 -209 259 -195
rect 280 -200 284 -195
rect 274 -204 280 -200
rect 284 -204 290 -200
rect 280 -209 284 -204
rect 305 -209 308 -195
rect 256 -213 257 -209
rect 307 -213 308 -209
rect 256 -263 259 -213
rect 269 -223 272 -213
rect 292 -216 295 -213
rect 279 -219 295 -216
rect 269 -226 285 -223
rect 269 -228 272 -226
rect 292 -228 295 -219
rect 280 -236 284 -233
rect 272 -240 280 -236
rect 284 -240 292 -236
rect 280 -243 284 -240
rect 269 -250 272 -248
rect 269 -253 285 -250
rect 269 -263 272 -253
rect 292 -257 295 -248
rect 279 -260 295 -257
rect 292 -263 295 -260
rect 305 -263 308 -213
rect 256 -267 257 -263
rect 307 -267 308 -263
rect 256 -281 259 -267
rect 280 -272 284 -267
rect 274 -276 280 -272
rect 284 -276 290 -272
rect 280 -281 284 -276
rect 305 -281 308 -267
rect 256 -285 257 -281
rect 307 -285 308 -281
rect 256 -335 259 -285
rect 269 -295 272 -285
rect 292 -288 295 -285
rect 279 -291 295 -288
rect 269 -298 285 -295
rect 269 -300 272 -298
rect 292 -300 295 -291
rect 280 -308 284 -305
rect 272 -312 280 -308
rect 284 -312 292 -308
rect 280 -315 284 -312
rect 269 -322 272 -320
rect 269 -325 285 -322
rect 269 -335 272 -325
rect 292 -329 295 -320
rect 279 -332 295 -329
rect 292 -335 295 -332
rect 305 -335 308 -285
rect 256 -339 257 -335
rect 307 -339 308 -335
rect 256 -353 259 -339
rect 280 -344 284 -339
rect 274 -348 280 -344
rect 284 -348 290 -344
rect 280 -353 284 -348
rect 305 -353 308 -339
rect 256 -357 257 -353
rect 307 -357 308 -353
rect 256 -387 259 -357
rect 269 -367 272 -357
rect 292 -360 295 -357
rect 279 -363 295 -360
rect 269 -370 285 -367
rect 269 -372 272 -370
rect 292 -372 295 -363
rect 280 -380 284 -377
rect 272 -384 280 -380
rect 284 -384 292 -380
rect 305 -387 308 -357
rect 311 -119 314 -92
rect 327 -96 335 -92
rect 339 -96 347 -92
rect 335 -99 339 -96
rect 324 -106 327 -104
rect 324 -109 340 -106
rect 324 -119 327 -109
rect 347 -113 350 -104
rect 334 -116 350 -113
rect 347 -119 350 -116
rect 360 -119 363 -92
rect 311 -123 312 -119
rect 362 -123 363 -119
rect 311 -137 314 -123
rect 335 -128 339 -123
rect 329 -132 335 -128
rect 339 -132 345 -128
rect 335 -137 339 -132
rect 360 -137 363 -123
rect 311 -141 312 -137
rect 362 -141 363 -137
rect 311 -191 314 -141
rect 324 -151 327 -141
rect 347 -144 350 -141
rect 334 -147 350 -144
rect 324 -154 340 -151
rect 324 -156 327 -154
rect 347 -156 350 -147
rect 335 -164 339 -161
rect 327 -168 335 -164
rect 339 -168 347 -164
rect 335 -171 339 -168
rect 324 -178 327 -176
rect 324 -181 340 -178
rect 324 -191 327 -181
rect 347 -185 350 -176
rect 334 -188 350 -185
rect 347 -191 350 -188
rect 360 -191 363 -141
rect 311 -195 312 -191
rect 362 -195 363 -191
rect 311 -209 314 -195
rect 335 -200 339 -195
rect 329 -204 335 -200
rect 339 -204 345 -200
rect 335 -209 339 -204
rect 360 -209 363 -195
rect 311 -213 312 -209
rect 362 -213 363 -209
rect 311 -263 314 -213
rect 324 -223 327 -213
rect 347 -216 350 -213
rect 334 -219 350 -216
rect 324 -226 340 -223
rect 324 -228 327 -226
rect 347 -228 350 -219
rect 335 -236 339 -233
rect 327 -240 335 -236
rect 339 -240 347 -236
rect 335 -243 339 -240
rect 324 -250 327 -248
rect 324 -253 340 -250
rect 324 -263 327 -253
rect 347 -257 350 -248
rect 334 -260 350 -257
rect 347 -263 350 -260
rect 360 -263 363 -213
rect 311 -267 312 -263
rect 362 -267 363 -263
rect 311 -281 314 -267
rect 335 -272 339 -267
rect 329 -276 335 -272
rect 339 -276 345 -272
rect 335 -281 339 -276
rect 360 -281 363 -267
rect 311 -285 312 -281
rect 362 -285 363 -281
rect 311 -335 314 -285
rect 324 -295 327 -285
rect 347 -288 350 -285
rect 334 -291 350 -288
rect 324 -298 340 -295
rect 324 -300 327 -298
rect 347 -300 350 -291
rect 335 -308 339 -305
rect 327 -312 335 -308
rect 339 -312 347 -308
rect 335 -315 339 -312
rect 324 -322 327 -320
rect 324 -325 340 -322
rect 324 -335 327 -325
rect 347 -329 350 -320
rect 334 -332 350 -329
rect 347 -335 350 -332
rect 360 -335 363 -285
rect 311 -339 312 -335
rect 362 -339 363 -335
rect 311 -353 314 -339
rect 335 -344 339 -339
rect 329 -348 335 -344
rect 339 -348 345 -344
rect 335 -353 339 -348
rect 360 -353 363 -339
rect 311 -357 312 -353
rect 362 -357 363 -353
rect 311 -387 314 -357
rect 324 -367 327 -357
rect 347 -360 350 -357
rect 334 -363 350 -360
rect 324 -370 340 -367
rect 324 -372 327 -370
rect 347 -372 350 -363
rect 335 -380 339 -377
rect 327 -384 335 -380
rect 339 -384 347 -380
rect 360 -387 363 -357
rect 366 -119 369 -92
rect 382 -96 390 -92
rect 394 -96 402 -92
rect 390 -99 394 -96
rect 379 -106 382 -104
rect 379 -109 395 -106
rect 379 -119 382 -109
rect 402 -113 405 -104
rect 389 -116 405 -113
rect 402 -119 405 -116
rect 415 -119 418 -92
rect 366 -123 367 -119
rect 417 -123 418 -119
rect 366 -137 369 -123
rect 390 -128 394 -123
rect 384 -132 390 -128
rect 394 -132 400 -128
rect 390 -137 394 -132
rect 415 -137 418 -123
rect 366 -141 367 -137
rect 417 -141 418 -137
rect 366 -191 369 -141
rect 379 -151 382 -141
rect 402 -144 405 -141
rect 389 -147 405 -144
rect 379 -154 395 -151
rect 379 -156 382 -154
rect 402 -156 405 -147
rect 390 -164 394 -161
rect 382 -168 390 -164
rect 394 -168 402 -164
rect 390 -171 394 -168
rect 379 -178 382 -176
rect 379 -181 395 -178
rect 379 -191 382 -181
rect 402 -185 405 -176
rect 389 -188 405 -185
rect 402 -191 405 -188
rect 415 -191 418 -141
rect 366 -195 367 -191
rect 417 -195 418 -191
rect 366 -209 369 -195
rect 390 -200 394 -195
rect 384 -204 390 -200
rect 394 -204 400 -200
rect 390 -209 394 -204
rect 415 -209 418 -195
rect 366 -213 367 -209
rect 417 -213 418 -209
rect 366 -263 369 -213
rect 379 -223 382 -213
rect 402 -216 405 -213
rect 389 -219 405 -216
rect 379 -226 395 -223
rect 379 -228 382 -226
rect 402 -228 405 -219
rect 390 -236 394 -233
rect 382 -240 390 -236
rect 394 -240 402 -236
rect 390 -243 394 -240
rect 379 -250 382 -248
rect 379 -253 395 -250
rect 379 -263 382 -253
rect 402 -257 405 -248
rect 389 -260 405 -257
rect 402 -263 405 -260
rect 415 -263 418 -213
rect 366 -267 367 -263
rect 417 -267 418 -263
rect 366 -281 369 -267
rect 390 -272 394 -267
rect 384 -276 390 -272
rect 394 -276 400 -272
rect 390 -281 394 -276
rect 415 -281 418 -267
rect 366 -285 367 -281
rect 417 -285 418 -281
rect 366 -335 369 -285
rect 379 -295 382 -285
rect 402 -288 405 -285
rect 389 -291 405 -288
rect 379 -298 395 -295
rect 379 -300 382 -298
rect 402 -300 405 -291
rect 390 -308 394 -305
rect 382 -312 390 -308
rect 394 -312 402 -308
rect 390 -315 394 -312
rect 379 -322 382 -320
rect 379 -325 395 -322
rect 379 -335 382 -325
rect 402 -329 405 -320
rect 389 -332 405 -329
rect 402 -335 405 -332
rect 415 -335 418 -285
rect 366 -339 367 -335
rect 417 -339 418 -335
rect 366 -353 369 -339
rect 390 -344 394 -339
rect 384 -348 390 -344
rect 394 -348 400 -344
rect 390 -353 394 -348
rect 415 -353 418 -339
rect 366 -357 367 -353
rect 417 -357 418 -353
rect 366 -387 369 -357
rect 379 -367 382 -357
rect 402 -360 405 -357
rect 389 -363 405 -360
rect 379 -370 395 -367
rect 379 -372 382 -370
rect 402 -372 405 -363
rect 390 -380 394 -377
rect 382 -384 390 -380
rect 394 -384 402 -380
rect 415 -387 418 -357
rect 421 -119 424 -92
rect 437 -96 445 -92
rect 449 -96 457 -92
rect 445 -99 449 -96
rect 434 -106 437 -104
rect 434 -109 450 -106
rect 434 -119 437 -109
rect 457 -113 460 -104
rect 444 -116 460 -113
rect 457 -119 460 -116
rect 470 -119 473 -92
rect 421 -123 422 -119
rect 472 -123 473 -119
rect 421 -137 424 -123
rect 445 -128 449 -123
rect 439 -132 445 -128
rect 449 -132 455 -128
rect 445 -137 449 -132
rect 470 -137 473 -123
rect 421 -141 422 -137
rect 472 -141 473 -137
rect 421 -191 424 -141
rect 434 -151 437 -141
rect 457 -144 460 -141
rect 444 -147 460 -144
rect 434 -154 450 -151
rect 434 -156 437 -154
rect 457 -156 460 -147
rect 445 -164 449 -161
rect 437 -168 445 -164
rect 449 -168 457 -164
rect 445 -171 449 -168
rect 434 -178 437 -176
rect 434 -181 450 -178
rect 434 -191 437 -181
rect 457 -185 460 -176
rect 444 -188 460 -185
rect 457 -191 460 -188
rect 470 -191 473 -141
rect 421 -195 422 -191
rect 472 -195 473 -191
rect 421 -209 424 -195
rect 445 -200 449 -195
rect 439 -204 445 -200
rect 449 -204 455 -200
rect 445 -209 449 -204
rect 470 -209 473 -195
rect 421 -213 422 -209
rect 472 -213 473 -209
rect 421 -263 424 -213
rect 434 -223 437 -213
rect 457 -216 460 -213
rect 444 -219 460 -216
rect 434 -226 450 -223
rect 434 -228 437 -226
rect 457 -228 460 -219
rect 445 -236 449 -233
rect 437 -240 445 -236
rect 449 -240 457 -236
rect 445 -243 449 -240
rect 434 -250 437 -248
rect 434 -253 450 -250
rect 434 -263 437 -253
rect 457 -257 460 -248
rect 444 -260 460 -257
rect 457 -263 460 -260
rect 470 -263 473 -213
rect 421 -267 422 -263
rect 472 -267 473 -263
rect 421 -281 424 -267
rect 445 -272 449 -267
rect 439 -276 445 -272
rect 449 -276 455 -272
rect 445 -281 449 -276
rect 470 -281 473 -267
rect 421 -285 422 -281
rect 472 -285 473 -281
rect 421 -335 424 -285
rect 434 -295 437 -285
rect 457 -288 460 -285
rect 444 -291 460 -288
rect 434 -298 450 -295
rect 434 -300 437 -298
rect 457 -300 460 -291
rect 445 -308 449 -305
rect 437 -312 445 -308
rect 449 -312 457 -308
rect 445 -315 449 -312
rect 434 -322 437 -320
rect 434 -325 450 -322
rect 434 -335 437 -325
rect 457 -329 460 -320
rect 444 -332 460 -329
rect 457 -335 460 -332
rect 470 -335 473 -285
rect 421 -339 422 -335
rect 472 -339 473 -335
rect 421 -353 424 -339
rect 445 -344 449 -339
rect 439 -348 445 -344
rect 449 -348 455 -344
rect 445 -353 449 -348
rect 470 -353 473 -339
rect 421 -357 422 -353
rect 472 -357 473 -353
rect 421 -387 424 -357
rect 434 -367 437 -357
rect 457 -360 460 -357
rect 444 -363 460 -360
rect 434 -370 450 -367
rect 434 -372 437 -370
rect 457 -372 460 -363
rect 445 -380 449 -377
rect 437 -384 445 -380
rect 449 -384 457 -380
rect 470 -387 473 -357
rect 476 -119 479 -92
rect 492 -96 500 -92
rect 504 -96 512 -92
rect 500 -99 504 -96
rect 489 -106 492 -104
rect 489 -109 505 -106
rect 489 -119 492 -109
rect 512 -113 515 -104
rect 499 -116 515 -113
rect 512 -119 515 -116
rect 525 -119 528 -92
rect 476 -123 477 -119
rect 527 -123 528 -119
rect 476 -137 479 -123
rect 500 -128 504 -123
rect 494 -132 500 -128
rect 504 -132 510 -128
rect 500 -137 504 -132
rect 525 -137 528 -123
rect 476 -141 477 -137
rect 527 -141 528 -137
rect 476 -191 479 -141
rect 489 -151 492 -141
rect 512 -144 515 -141
rect 499 -147 515 -144
rect 489 -154 505 -151
rect 489 -156 492 -154
rect 512 -156 515 -147
rect 500 -164 504 -161
rect 492 -168 500 -164
rect 504 -168 512 -164
rect 500 -171 504 -168
rect 489 -178 492 -176
rect 489 -181 505 -178
rect 489 -191 492 -181
rect 512 -185 515 -176
rect 499 -188 515 -185
rect 512 -191 515 -188
rect 525 -191 528 -141
rect 476 -195 477 -191
rect 527 -195 528 -191
rect 476 -209 479 -195
rect 500 -200 504 -195
rect 494 -204 500 -200
rect 504 -204 510 -200
rect 500 -209 504 -204
rect 525 -209 528 -195
rect 476 -213 477 -209
rect 527 -213 528 -209
rect 476 -263 479 -213
rect 489 -223 492 -213
rect 512 -216 515 -213
rect 499 -219 515 -216
rect 489 -226 505 -223
rect 489 -228 492 -226
rect 512 -228 515 -219
rect 500 -236 504 -233
rect 492 -240 500 -236
rect 504 -240 512 -236
rect 500 -243 504 -240
rect 489 -250 492 -248
rect 489 -253 505 -250
rect 489 -263 492 -253
rect 512 -257 515 -248
rect 499 -260 515 -257
rect 512 -263 515 -260
rect 525 -263 528 -213
rect 476 -267 477 -263
rect 527 -267 528 -263
rect 476 -281 479 -267
rect 500 -272 504 -267
rect 494 -276 500 -272
rect 504 -276 510 -272
rect 500 -281 504 -276
rect 525 -281 528 -267
rect 476 -285 477 -281
rect 527 -285 528 -281
rect 476 -335 479 -285
rect 489 -295 492 -285
rect 512 -288 515 -285
rect 499 -291 515 -288
rect 489 -298 505 -295
rect 489 -300 492 -298
rect 512 -300 515 -291
rect 500 -308 504 -305
rect 492 -312 500 -308
rect 504 -312 512 -308
rect 500 -315 504 -312
rect 489 -322 492 -320
rect 489 -325 505 -322
rect 489 -335 492 -325
rect 512 -329 515 -320
rect 499 -332 515 -329
rect 512 -335 515 -332
rect 525 -335 528 -285
rect 476 -339 477 -335
rect 527 -339 528 -335
rect 476 -353 479 -339
rect 500 -344 504 -339
rect 494 -348 500 -344
rect 504 -348 510 -344
rect 500 -353 504 -348
rect 525 -353 528 -339
rect 476 -357 477 -353
rect 527 -357 528 -353
rect 476 -387 479 -357
rect 489 -367 492 -357
rect 512 -360 515 -357
rect 499 -363 515 -360
rect 489 -370 505 -367
rect 489 -372 492 -370
rect 512 -372 515 -363
rect 500 -380 504 -377
rect 492 -384 500 -380
rect 504 -384 512 -380
rect 525 -387 528 -357
rect 531 -119 534 -92
rect 547 -96 555 -92
rect 559 -96 567 -92
rect 555 -99 559 -96
rect 544 -106 547 -104
rect 544 -109 560 -106
rect 544 -119 547 -109
rect 567 -113 570 -104
rect 554 -116 570 -113
rect 567 -119 570 -116
rect 580 -119 583 -92
rect 531 -123 532 -119
rect 582 -123 583 -119
rect 531 -137 534 -123
rect 555 -128 559 -123
rect 549 -132 555 -128
rect 559 -132 565 -128
rect 555 -137 559 -132
rect 580 -137 583 -123
rect 531 -141 532 -137
rect 582 -141 583 -137
rect 531 -191 534 -141
rect 544 -151 547 -141
rect 567 -144 570 -141
rect 554 -147 570 -144
rect 544 -154 560 -151
rect 544 -156 547 -154
rect 567 -156 570 -147
rect 555 -164 559 -161
rect 547 -168 555 -164
rect 559 -168 567 -164
rect 555 -171 559 -168
rect 544 -178 547 -176
rect 544 -181 560 -178
rect 544 -191 547 -181
rect 567 -185 570 -176
rect 554 -188 570 -185
rect 567 -191 570 -188
rect 580 -191 583 -141
rect 531 -195 532 -191
rect 582 -195 583 -191
rect 531 -209 534 -195
rect 555 -200 559 -195
rect 549 -204 555 -200
rect 559 -204 565 -200
rect 555 -209 559 -204
rect 580 -209 583 -195
rect 531 -213 532 -209
rect 582 -213 583 -209
rect 531 -263 534 -213
rect 544 -223 547 -213
rect 567 -216 570 -213
rect 554 -219 570 -216
rect 544 -226 560 -223
rect 544 -228 547 -226
rect 567 -228 570 -219
rect 555 -236 559 -233
rect 547 -240 555 -236
rect 559 -240 567 -236
rect 555 -243 559 -240
rect 544 -250 547 -248
rect 544 -253 560 -250
rect 544 -263 547 -253
rect 567 -257 570 -248
rect 554 -260 570 -257
rect 567 -263 570 -260
rect 580 -263 583 -213
rect 531 -267 532 -263
rect 582 -267 583 -263
rect 531 -281 534 -267
rect 555 -272 559 -267
rect 549 -276 555 -272
rect 559 -276 565 -272
rect 555 -281 559 -276
rect 580 -281 583 -267
rect 531 -285 532 -281
rect 582 -285 583 -281
rect 531 -335 534 -285
rect 544 -295 547 -285
rect 567 -288 570 -285
rect 554 -291 570 -288
rect 544 -298 560 -295
rect 544 -300 547 -298
rect 567 -300 570 -291
rect 555 -308 559 -305
rect 547 -312 555 -308
rect 559 -312 567 -308
rect 555 -315 559 -312
rect 544 -322 547 -320
rect 544 -325 560 -322
rect 544 -335 547 -325
rect 567 -329 570 -320
rect 554 -332 570 -329
rect 567 -335 570 -332
rect 580 -335 583 -285
rect 531 -339 532 -335
rect 582 -339 583 -335
rect 531 -353 534 -339
rect 555 -344 559 -339
rect 549 -348 555 -344
rect 559 -348 565 -344
rect 555 -353 559 -348
rect 580 -353 583 -339
rect 531 -357 532 -353
rect 582 -357 583 -353
rect 531 -387 534 -357
rect 544 -367 547 -357
rect 567 -360 570 -357
rect 554 -363 570 -360
rect 544 -370 560 -367
rect 544 -372 547 -370
rect 567 -372 570 -363
rect 555 -380 559 -377
rect 547 -384 555 -380
rect 559 -384 567 -380
rect 580 -387 583 -357
rect 586 -119 589 -92
rect 602 -96 610 -92
rect 614 -96 622 -92
rect 610 -99 614 -96
rect 599 -106 602 -104
rect 599 -109 615 -106
rect 599 -119 602 -109
rect 622 -113 625 -104
rect 609 -116 625 -113
rect 622 -119 625 -116
rect 635 -119 638 -92
rect 586 -123 587 -119
rect 637 -123 638 -119
rect 586 -137 589 -123
rect 610 -128 614 -123
rect 604 -132 610 -128
rect 614 -132 620 -128
rect 610 -137 614 -132
rect 635 -137 638 -123
rect 586 -141 587 -137
rect 637 -141 638 -137
rect 586 -191 589 -141
rect 599 -151 602 -141
rect 622 -144 625 -141
rect 609 -147 625 -144
rect 599 -154 615 -151
rect 599 -156 602 -154
rect 622 -156 625 -147
rect 610 -164 614 -161
rect 602 -168 610 -164
rect 614 -168 622 -164
rect 610 -171 614 -168
rect 599 -178 602 -176
rect 599 -181 615 -178
rect 599 -191 602 -181
rect 622 -185 625 -176
rect 609 -188 625 -185
rect 622 -191 625 -188
rect 635 -191 638 -141
rect 586 -195 587 -191
rect 637 -195 638 -191
rect 586 -209 589 -195
rect 610 -200 614 -195
rect 604 -204 610 -200
rect 614 -204 620 -200
rect 610 -209 614 -204
rect 635 -209 638 -195
rect 586 -213 587 -209
rect 637 -213 638 -209
rect 586 -263 589 -213
rect 599 -223 602 -213
rect 622 -216 625 -213
rect 609 -219 625 -216
rect 599 -226 615 -223
rect 599 -228 602 -226
rect 622 -228 625 -219
rect 610 -236 614 -233
rect 602 -240 610 -236
rect 614 -240 622 -236
rect 610 -243 614 -240
rect 599 -250 602 -248
rect 599 -253 615 -250
rect 599 -263 602 -253
rect 622 -257 625 -248
rect 609 -260 625 -257
rect 622 -263 625 -260
rect 635 -263 638 -213
rect 586 -267 587 -263
rect 637 -267 638 -263
rect 586 -281 589 -267
rect 610 -272 614 -267
rect 604 -276 610 -272
rect 614 -276 620 -272
rect 610 -281 614 -276
rect 635 -281 638 -267
rect 586 -285 587 -281
rect 637 -285 638 -281
rect 586 -335 589 -285
rect 599 -295 602 -285
rect 622 -288 625 -285
rect 609 -291 625 -288
rect 599 -298 615 -295
rect 599 -300 602 -298
rect 622 -300 625 -291
rect 610 -308 614 -305
rect 602 -312 610 -308
rect 614 -312 622 -308
rect 610 -315 614 -312
rect 599 -322 602 -320
rect 599 -325 615 -322
rect 599 -335 602 -325
rect 622 -329 625 -320
rect 609 -332 625 -329
rect 622 -335 625 -332
rect 635 -335 638 -285
rect 586 -339 587 -335
rect 637 -339 638 -335
rect 586 -353 589 -339
rect 610 -344 614 -339
rect 604 -348 610 -344
rect 614 -348 620 -344
rect 610 -353 614 -348
rect 635 -353 638 -339
rect 586 -357 587 -353
rect 637 -357 638 -353
rect 586 -387 589 -357
rect 599 -367 602 -357
rect 622 -360 625 -357
rect 609 -363 625 -360
rect 599 -370 615 -367
rect 599 -372 602 -370
rect 622 -372 625 -363
rect 610 -380 614 -377
rect 602 -384 610 -380
rect 614 -384 622 -380
rect 635 -387 638 -357
<< m2contact >>
rect 225 -96 229 -92
rect 207 -114 211 -110
rect 243 -114 247 -110
rect 225 -132 229 -128
rect 207 -150 211 -146
rect 243 -150 247 -146
rect 225 -168 229 -164
rect 207 -186 211 -182
rect 243 -186 247 -182
rect 225 -204 229 -200
rect 207 -222 211 -218
rect 243 -222 247 -218
rect 225 -240 229 -236
rect 207 -258 211 -254
rect 243 -258 247 -254
rect 225 -276 229 -272
rect 207 -294 211 -290
rect 243 -294 247 -290
rect 225 -312 229 -308
rect 207 -330 211 -326
rect 243 -330 247 -326
rect 225 -348 229 -344
rect 207 -366 211 -362
rect 243 -366 247 -362
rect 225 -384 229 -380
rect 280 -96 284 -92
rect 262 -114 266 -110
rect 298 -114 302 -110
rect 280 -132 284 -128
rect 262 -150 266 -146
rect 298 -150 302 -146
rect 280 -168 284 -164
rect 262 -186 266 -182
rect 298 -186 302 -182
rect 280 -204 284 -200
rect 262 -222 266 -218
rect 298 -222 302 -218
rect 280 -240 284 -236
rect 262 -258 266 -254
rect 298 -258 302 -254
rect 280 -276 284 -272
rect 262 -294 266 -290
rect 298 -294 302 -290
rect 280 -312 284 -308
rect 262 -330 266 -326
rect 298 -330 302 -326
rect 280 -348 284 -344
rect 262 -366 266 -362
rect 298 -366 302 -362
rect 280 -384 284 -380
rect 335 -96 339 -92
rect 317 -114 321 -110
rect 353 -114 357 -110
rect 335 -132 339 -128
rect 317 -150 321 -146
rect 353 -150 357 -146
rect 335 -168 339 -164
rect 317 -186 321 -182
rect 353 -186 357 -182
rect 335 -204 339 -200
rect 317 -222 321 -218
rect 353 -222 357 -218
rect 335 -240 339 -236
rect 317 -258 321 -254
rect 353 -258 357 -254
rect 335 -276 339 -272
rect 317 -294 321 -290
rect 353 -294 357 -290
rect 335 -312 339 -308
rect 317 -330 321 -326
rect 353 -330 357 -326
rect 335 -348 339 -344
rect 317 -366 321 -362
rect 353 -366 357 -362
rect 335 -384 339 -380
rect 390 -96 394 -92
rect 372 -114 376 -110
rect 408 -114 412 -110
rect 390 -132 394 -128
rect 372 -150 376 -146
rect 408 -150 412 -146
rect 390 -168 394 -164
rect 372 -186 376 -182
rect 408 -186 412 -182
rect 390 -204 394 -200
rect 372 -222 376 -218
rect 408 -222 412 -218
rect 390 -240 394 -236
rect 372 -258 376 -254
rect 408 -258 412 -254
rect 390 -276 394 -272
rect 372 -294 376 -290
rect 408 -294 412 -290
rect 390 -312 394 -308
rect 372 -330 376 -326
rect 408 -330 412 -326
rect 390 -348 394 -344
rect 372 -366 376 -362
rect 408 -366 412 -362
rect 390 -384 394 -380
rect 445 -96 449 -92
rect 427 -114 431 -110
rect 463 -114 467 -110
rect 445 -132 449 -128
rect 427 -150 431 -146
rect 463 -150 467 -146
rect 445 -168 449 -164
rect 427 -186 431 -182
rect 463 -186 467 -182
rect 445 -204 449 -200
rect 427 -222 431 -218
rect 463 -222 467 -218
rect 445 -240 449 -236
rect 427 -258 431 -254
rect 463 -258 467 -254
rect 445 -276 449 -272
rect 427 -294 431 -290
rect 463 -294 467 -290
rect 445 -312 449 -308
rect 427 -330 431 -326
rect 463 -330 467 -326
rect 445 -348 449 -344
rect 427 -366 431 -362
rect 463 -366 467 -362
rect 445 -384 449 -380
rect 500 -96 504 -92
rect 482 -114 486 -110
rect 518 -114 522 -110
rect 500 -132 504 -128
rect 482 -150 486 -146
rect 518 -150 522 -146
rect 500 -168 504 -164
rect 482 -186 486 -182
rect 518 -186 522 -182
rect 500 -204 504 -200
rect 482 -222 486 -218
rect 518 -222 522 -218
rect 500 -240 504 -236
rect 482 -258 486 -254
rect 518 -258 522 -254
rect 500 -276 504 -272
rect 482 -294 486 -290
rect 518 -294 522 -290
rect 500 -312 504 -308
rect 482 -330 486 -326
rect 518 -330 522 -326
rect 500 -348 504 -344
rect 482 -366 486 -362
rect 518 -366 522 -362
rect 500 -384 504 -380
rect 555 -96 559 -92
rect 537 -114 541 -110
rect 573 -114 577 -110
rect 555 -132 559 -128
rect 537 -150 541 -146
rect 573 -150 577 -146
rect 555 -168 559 -164
rect 537 -186 541 -182
rect 573 -186 577 -182
rect 555 -204 559 -200
rect 537 -222 541 -218
rect 573 -222 577 -218
rect 555 -240 559 -236
rect 537 -258 541 -254
rect 573 -258 577 -254
rect 555 -276 559 -272
rect 537 -294 541 -290
rect 573 -294 577 -290
rect 555 -312 559 -308
rect 537 -330 541 -326
rect 573 -330 577 -326
rect 555 -348 559 -344
rect 537 -366 541 -362
rect 573 -366 577 -362
rect 555 -384 559 -380
rect 610 -96 614 -92
rect 592 -114 596 -110
rect 628 -114 632 -110
rect 610 -132 614 -128
rect 592 -150 596 -146
rect 628 -150 632 -146
rect 610 -168 614 -164
rect 592 -186 596 -182
rect 628 -186 632 -182
rect 610 -204 614 -200
rect 592 -222 596 -218
rect 628 -222 632 -218
rect 610 -240 614 -236
rect 592 -258 596 -254
rect 628 -258 632 -254
rect 610 -276 614 -272
rect 592 -294 596 -290
rect 628 -294 632 -290
rect 610 -312 614 -308
rect 592 -330 596 -326
rect 628 -330 632 -326
rect 610 -348 614 -344
rect 592 -366 596 -362
rect 628 -366 632 -362
rect 610 -384 614 -380
<< metal2 >>
rect 198 -96 225 -92
rect 229 -96 280 -92
rect 284 -96 335 -92
rect 339 -96 390 -92
rect 394 -96 445 -92
rect 449 -96 500 -92
rect 504 -96 555 -92
rect 559 -96 610 -92
rect 614 -96 641 -92
rect 198 -114 207 -110
rect 211 -114 243 -110
rect 247 -114 262 -110
rect 266 -114 298 -110
rect 302 -114 317 -110
rect 321 -114 353 -110
rect 357 -114 372 -110
rect 376 -114 408 -110
rect 412 -114 427 -110
rect 431 -114 463 -110
rect 467 -114 482 -110
rect 486 -114 518 -110
rect 522 -114 537 -110
rect 541 -114 573 -110
rect 577 -114 592 -110
rect 596 -114 628 -110
rect 632 -114 641 -110
rect 198 -132 225 -128
rect 229 -132 280 -128
rect 284 -132 335 -128
rect 339 -132 390 -128
rect 394 -132 445 -128
rect 449 -132 500 -128
rect 504 -132 555 -128
rect 559 -132 610 -128
rect 614 -132 641 -128
rect 198 -150 207 -146
rect 211 -150 243 -146
rect 247 -150 262 -146
rect 266 -150 298 -146
rect 302 -150 317 -146
rect 321 -150 353 -146
rect 357 -150 372 -146
rect 376 -150 408 -146
rect 412 -150 427 -146
rect 431 -150 463 -146
rect 467 -150 482 -146
rect 486 -150 518 -146
rect 522 -150 537 -146
rect 541 -150 573 -146
rect 577 -150 592 -146
rect 596 -150 628 -146
rect 632 -150 641 -146
rect 198 -168 225 -164
rect 229 -168 280 -164
rect 284 -168 335 -164
rect 339 -168 390 -164
rect 394 -168 445 -164
rect 449 -168 500 -164
rect 504 -168 555 -164
rect 559 -168 610 -164
rect 614 -168 641 -164
rect 198 -186 207 -182
rect 211 -186 243 -182
rect 247 -186 262 -182
rect 266 -186 298 -182
rect 302 -186 317 -182
rect 321 -186 353 -182
rect 357 -186 372 -182
rect 376 -186 408 -182
rect 412 -186 427 -182
rect 431 -186 463 -182
rect 467 -186 482 -182
rect 486 -186 518 -182
rect 522 -186 537 -182
rect 541 -186 573 -182
rect 577 -186 592 -182
rect 596 -186 628 -182
rect 632 -186 641 -182
rect 198 -204 225 -200
rect 229 -204 280 -200
rect 284 -204 335 -200
rect 339 -204 390 -200
rect 394 -204 445 -200
rect 449 -204 500 -200
rect 504 -204 555 -200
rect 559 -204 610 -200
rect 614 -204 641 -200
rect 198 -222 207 -218
rect 211 -222 243 -218
rect 247 -222 262 -218
rect 266 -222 298 -218
rect 302 -222 317 -218
rect 321 -222 353 -218
rect 357 -222 372 -218
rect 376 -222 408 -218
rect 412 -222 427 -218
rect 431 -222 463 -218
rect 467 -222 482 -218
rect 486 -222 518 -218
rect 522 -222 537 -218
rect 541 -222 573 -218
rect 577 -222 592 -218
rect 596 -222 628 -218
rect 632 -222 641 -218
rect 198 -240 225 -236
rect 229 -240 280 -236
rect 284 -240 335 -236
rect 339 -240 390 -236
rect 394 -240 445 -236
rect 449 -240 500 -236
rect 504 -240 555 -236
rect 559 -240 610 -236
rect 614 -240 641 -236
rect 198 -258 207 -254
rect 211 -258 243 -254
rect 247 -258 262 -254
rect 266 -258 298 -254
rect 302 -258 317 -254
rect 321 -258 353 -254
rect 357 -258 372 -254
rect 376 -258 408 -254
rect 412 -258 427 -254
rect 431 -258 463 -254
rect 467 -258 482 -254
rect 486 -258 518 -254
rect 522 -258 537 -254
rect 541 -258 573 -254
rect 577 -258 592 -254
rect 596 -258 628 -254
rect 632 -258 641 -254
rect 198 -276 225 -272
rect 229 -276 280 -272
rect 284 -276 335 -272
rect 339 -276 390 -272
rect 394 -276 445 -272
rect 449 -276 500 -272
rect 504 -276 555 -272
rect 559 -276 610 -272
rect 614 -276 641 -272
rect 198 -294 207 -290
rect 211 -294 243 -290
rect 247 -294 262 -290
rect 266 -294 298 -290
rect 302 -294 317 -290
rect 321 -294 353 -290
rect 357 -294 372 -290
rect 376 -294 408 -290
rect 412 -294 427 -290
rect 431 -294 463 -290
rect 467 -294 482 -290
rect 486 -294 518 -290
rect 522 -294 537 -290
rect 541 -294 573 -290
rect 577 -294 592 -290
rect 596 -294 628 -290
rect 632 -294 641 -290
rect 198 -312 225 -308
rect 229 -312 280 -308
rect 284 -312 335 -308
rect 339 -312 390 -308
rect 394 -312 445 -308
rect 449 -312 500 -308
rect 504 -312 555 -308
rect 559 -312 610 -308
rect 614 -312 641 -308
rect 198 -330 207 -326
rect 211 -330 243 -326
rect 247 -330 262 -326
rect 266 -330 298 -326
rect 302 -330 317 -326
rect 321 -330 353 -326
rect 357 -330 372 -326
rect 376 -330 408 -326
rect 412 -330 427 -326
rect 431 -330 463 -326
rect 467 -330 482 -326
rect 486 -330 518 -326
rect 522 -330 537 -326
rect 541 -330 573 -326
rect 577 -330 592 -326
rect 596 -330 628 -326
rect 632 -330 641 -326
rect 198 -348 225 -344
rect 229 -348 280 -344
rect 284 -348 335 -344
rect 339 -348 390 -344
rect 394 -348 445 -344
rect 449 -348 500 -344
rect 504 -348 555 -344
rect 559 -348 610 -344
rect 614 -348 641 -344
rect 198 -366 207 -362
rect 211 -366 243 -362
rect 247 -366 262 -362
rect 266 -366 298 -362
rect 302 -366 317 -362
rect 321 -366 353 -362
rect 357 -366 372 -362
rect 376 -366 408 -362
rect 412 -366 427 -362
rect 431 -366 463 -362
rect 467 -366 482 -362
rect 486 -366 518 -362
rect 522 -366 537 -362
rect 541 -366 573 -362
rect 577 -366 592 -362
rect 596 -366 628 -362
rect 632 -366 641 -362
rect 198 -384 225 -380
rect 229 -384 280 -380
rect 284 -384 335 -380
rect 339 -384 390 -380
rect 394 -384 445 -380
rect 449 -384 500 -380
rect 504 -384 555 -380
rect 559 -384 610 -380
rect 614 -384 641 -380
use wd  wd_1 ~/lab/magic/sram/wd
timestamp 1635738960
transform 1 0 340 0 1 -202
box -283 -50 -223 64
use wd  wd_0
timestamp 1635738960
transform 1 0 285 0 1 -202
box -283 -50 -223 64
use sa  sa_1 ~/lab/magic/sram/sa
timestamp 1635742126
transform 1 0 83 0 1 -4
box -25 -131 33 -62
use sa  sa_0
timestamp 1635742126
transform 1 0 28 0 1 -4
box -25 -131 33 -62
use 6T-cell  6T-cell_3 ~/lab/magic/sram/6T-cell
timestamp 1635593005
transform 1 0 11 0 -1 -33
box 47 -8 105 38
use 6T-cell  6T-cell_2
timestamp 1635593005
transform 1 0 11 0 1 -27
box 47 -8 105 38
use 6T-cell  6T-cell_1
timestamp 1635593005
transform 1 0 -44 0 -1 -33
box 47 -8 105 38
use 6T-cell  6T-cell_0
timestamp 1635593005
transform 1 0 -44 0 1 -27
box 47 -8 105 38
use pc  pc_1 ~/lab/magic/sram/pc
timestamp 1635740445
transform 1 0 58 0 1 51
box 0 -47 58 -8
use pc  pc_0
timestamp 1635740445
transform 1 0 3 0 1 51
box 0 -47 58 -8
<< labels >>
rlabel metal1 202 -228 203 -227 3 bl
rlabel metal1 251 -228 252 -227 7 blb
rlabel metal2 199 -220 199 -220 3 wl
rlabel metal1 215 -225 216 -224 5 q1
rlabel metal1 238 -225 239 -224 5 q2
rlabel m2contact 227 -202 227 -202 1 gnd
rlabel metal1 202 -177 203 -176 3 bl
rlabel metal1 251 -177 252 -176 7 blb
rlabel metal2 199 -184 199 -184 3 wl
rlabel metal1 215 -180 216 -179 1 q1
rlabel metal1 238 -180 239 -179 1 q2
rlabel metal1 312 -228 313 -227 3 bl
rlabel metal1 361 -228 362 -227 7 blb
rlabel metal2 309 -220 309 -220 3 wl
rlabel metal1 325 -225 326 -224 5 q1
rlabel metal1 348 -225 349 -224 5 q2
rlabel m2contact 337 -202 337 -202 1 gnd
rlabel metal1 312 -177 313 -176 3 bl
rlabel metal1 361 -177 362 -176 7 blb
rlabel metal2 309 -184 309 -184 3 wl
rlabel metal1 325 -180 326 -179 1 q1
rlabel metal1 348 -180 349 -179 1 q2
rlabel metal1 257 -177 258 -176 3 bl
rlabel metal1 306 -177 307 -176 7 blb
rlabel metal2 254 -184 254 -184 3 wl
rlabel metal1 270 -180 271 -179 1 q1
rlabel metal1 293 -180 294 -179 1 q2
rlabel metal1 422 -228 423 -227 3 bl
rlabel metal1 471 -228 472 -227 7 blb
rlabel metal2 419 -220 419 -220 3 wl
rlabel metal1 435 -225 436 -224 5 q1
rlabel metal1 458 -225 459 -224 5 q2
rlabel metal1 367 -228 368 -227 3 bl
rlabel metal1 416 -228 417 -227 7 blb
rlabel metal2 364 -220 364 -220 3 wl
rlabel metal1 380 -225 381 -224 5 q1
rlabel metal1 403 -225 404 -224 5 q2
rlabel m2contact 447 -202 447 -202 1 gnd
rlabel metal1 422 -177 423 -176 3 bl
rlabel metal1 471 -177 472 -176 7 blb
rlabel metal2 419 -184 419 -184 3 wl
rlabel metal1 435 -180 436 -179 1 q1
rlabel metal1 458 -180 459 -179 1 q2
rlabel m2contact 392 -202 392 -202 1 gnd
rlabel metal1 367 -177 368 -176 3 bl
rlabel metal1 416 -177 417 -176 7 blb
rlabel metal2 364 -184 364 -184 3 wl
rlabel metal1 380 -180 381 -179 1 q1
rlabel metal1 403 -180 404 -179 1 q2
rlabel metal1 587 -228 588 -227 3 bl
rlabel metal1 636 -228 637 -227 7 blb
rlabel metal2 584 -220 584 -220 3 wl
rlabel metal1 600 -225 601 -224 5 q1
rlabel metal1 623 -225 624 -224 5 q2
rlabel metal1 532 -228 533 -227 3 bl
rlabel metal1 581 -228 582 -227 7 blb
rlabel metal2 529 -220 529 -220 3 wl
rlabel metal1 545 -225 546 -224 5 q1
rlabel metal1 568 -225 569 -224 5 q2
rlabel metal1 477 -228 478 -227 3 bl
rlabel metal1 526 -228 527 -227 7 blb
rlabel metal2 474 -220 474 -220 3 wl
rlabel metal1 490 -225 491 -224 5 q1
rlabel metal1 513 -225 514 -224 5 q2
rlabel m2contact 612 -202 612 -202 1 gnd
rlabel metal1 587 -177 588 -176 3 bl
rlabel metal1 636 -177 637 -176 7 blb
rlabel metal2 584 -184 584 -184 3 wl
rlabel metal1 600 -180 601 -179 1 q1
rlabel metal1 623 -180 624 -179 1 q2
rlabel m2contact 557 -202 557 -202 1 gnd
rlabel metal1 532 -177 533 -176 3 bl
rlabel metal1 581 -177 582 -176 7 blb
rlabel metal2 529 -184 529 -184 3 wl
rlabel metal1 545 -180 546 -179 1 q1
rlabel metal1 568 -180 569 -179 1 q2
rlabel m2contact 502 -202 502 -202 1 gnd
rlabel metal1 477 -177 478 -176 3 bl
rlabel metal1 526 -177 527 -176 7 blb
rlabel metal2 474 -184 474 -184 3 wl
rlabel metal1 490 -180 491 -179 1 q1
rlabel metal1 513 -180 514 -179 1 q2
rlabel m2contact 282 -202 282 -202 5 gnd
rlabel metal1 257 -228 258 -227 3 bl
rlabel metal1 306 -228 307 -227 7 blb
rlabel metal2 254 -220 254 -220 3 wl
rlabel metal1 270 -225 271 -224 5 q1
rlabel metal1 293 -225 294 -224 5 q2
rlabel m2contact 227 -166 227 -166 1 vdd
rlabel metal1 202 -156 203 -155 3 bl
rlabel metal1 251 -156 252 -155 7 blb
rlabel metal2 199 -148 199 -148 3 wl
rlabel metal1 215 -153 216 -152 5 q1
rlabel metal1 238 -153 239 -152 5 q2
rlabel m2contact 337 -166 337 -166 1 vdd
rlabel metal1 312 -156 313 -155 3 bl
rlabel metal1 361 -156 362 -155 7 blb
rlabel metal2 309 -148 309 -148 3 wl
rlabel metal1 325 -153 326 -152 5 q1
rlabel metal1 348 -153 349 -152 5 q2
rlabel m2contact 282 -166 282 -166 1 vdd
rlabel metal1 257 -156 258 -155 3 bl
rlabel metal1 306 -156 307 -155 7 blb
rlabel metal2 254 -148 254 -148 3 wl
rlabel metal1 270 -153 271 -152 5 q1
rlabel metal1 293 -153 294 -152 5 q2
rlabel m2contact 447 -166 447 -166 1 vdd
rlabel metal1 422 -156 423 -155 3 bl
rlabel metal1 471 -156 472 -155 7 blb
rlabel metal2 419 -148 419 -148 3 wl
rlabel metal1 435 -153 436 -152 5 q1
rlabel metal1 458 -153 459 -152 5 q2
rlabel m2contact 392 -166 392 -166 1 vdd
rlabel metal1 367 -156 368 -155 3 bl
rlabel metal1 416 -156 417 -155 7 blb
rlabel metal2 364 -148 364 -148 3 wl
rlabel metal1 380 -153 381 -152 5 q1
rlabel metal1 403 -153 404 -152 5 q2
rlabel m2contact 612 -166 612 -166 1 vdd
rlabel metal1 587 -156 588 -155 3 bl
rlabel metal1 636 -156 637 -155 7 blb
rlabel metal2 584 -148 584 -148 3 wl
rlabel metal1 600 -153 601 -152 5 q1
rlabel metal1 623 -153 624 -152 5 q2
rlabel m2contact 557 -166 557 -166 1 vdd
rlabel metal1 532 -156 533 -155 3 bl
rlabel metal1 581 -156 582 -155 7 blb
rlabel metal2 529 -148 529 -148 3 wl
rlabel metal1 545 -153 546 -152 5 q1
rlabel metal1 568 -153 569 -152 5 q2
rlabel m2contact 502 -166 502 -166 1 vdd
rlabel metal1 477 -156 478 -155 3 bl
rlabel metal1 526 -156 527 -155 7 blb
rlabel metal2 474 -148 474 -148 3 wl
rlabel metal1 490 -153 491 -152 5 q1
rlabel metal1 513 -153 514 -152 5 q2
rlabel m2contact 227 -130 227 -130 1 gnd
rlabel metal1 202 -105 203 -104 3 bl
rlabel metal1 251 -105 252 -104 7 blb
rlabel metal2 199 -112 199 -112 3 wl
rlabel metal1 215 -108 216 -107 1 q1
rlabel metal1 238 -108 239 -107 1 q2
rlabel m2contact 337 -130 337 -130 1 gnd
rlabel metal1 312 -105 313 -104 3 bl
rlabel metal1 361 -105 362 -104 7 blb
rlabel metal2 309 -112 309 -112 3 wl
rlabel metal1 325 -108 326 -107 1 q1
rlabel metal1 348 -108 349 -107 1 q2
rlabel metal1 257 -105 258 -104 3 bl
rlabel metal1 306 -105 307 -104 7 blb
rlabel metal2 254 -112 254 -112 3 wl
rlabel metal1 270 -108 271 -107 1 q1
rlabel metal1 293 -108 294 -107 1 q2
rlabel m2contact 447 -130 447 -130 1 gnd
rlabel metal1 422 -105 423 -104 3 bl
rlabel metal1 471 -105 472 -104 7 blb
rlabel metal2 419 -112 419 -112 3 wl
rlabel metal1 435 -108 436 -107 1 q1
rlabel metal1 458 -108 459 -107 1 q2
rlabel m2contact 392 -130 392 -130 1 gnd
rlabel metal1 367 -105 368 -104 3 bl
rlabel metal1 416 -105 417 -104 7 blb
rlabel metal2 364 -112 364 -112 3 wl
rlabel metal1 380 -108 381 -107 1 q1
rlabel metal1 403 -108 404 -107 1 q2
rlabel m2contact 612 -130 612 -130 1 gnd
rlabel metal1 587 -105 588 -104 3 bl
rlabel metal1 636 -105 637 -104 7 blb
rlabel metal2 584 -112 584 -112 3 wl
rlabel metal1 600 -108 601 -107 1 q1
rlabel metal1 623 -108 624 -107 1 q2
rlabel m2contact 557 -130 557 -130 1 gnd
rlabel metal1 532 -105 533 -104 3 bl
rlabel metal1 581 -105 582 -104 7 blb
rlabel metal2 529 -112 529 -112 3 wl
rlabel metal1 545 -108 546 -107 1 q1
rlabel metal1 568 -108 569 -107 1 q2
rlabel m2contact 502 -130 502 -130 1 gnd
rlabel metal1 477 -105 478 -104 3 bl
rlabel metal1 526 -105 527 -104 7 blb
rlabel metal2 474 -112 474 -112 3 wl
rlabel metal1 490 -108 491 -107 1 q1
rlabel metal1 513 -108 514 -107 1 q2
rlabel m2contact 282 -130 282 -130 5 gnd
rlabel m2contact 227 -94 227 -94 1 vdd
rlabel m2contact 337 -94 337 -94 1 vdd
rlabel m2contact 282 -94 282 -94 1 vdd
rlabel m2contact 447 -94 447 -94 1 vdd
rlabel m2contact 392 -94 392 -94 1 vdd
rlabel m2contact 612 -94 612 -94 1 vdd
rlabel m2contact 557 -94 557 -94 1 vdd
rlabel m2contact 502 -94 502 -94 1 vdd
rlabel m2contact 227 -382 227 -382 1 vdd
rlabel metal1 202 -372 203 -371 3 bl
rlabel metal1 251 -372 252 -371 7 blb
rlabel metal2 199 -364 199 -364 3 wl
rlabel metal1 215 -369 216 -368 5 q1
rlabel metal1 238 -369 239 -368 5 q2
rlabel m2contact 227 -346 227 -346 1 gnd
rlabel metal1 202 -321 203 -320 3 bl
rlabel metal1 251 -321 252 -320 7 blb
rlabel metal2 199 -328 199 -328 3 wl
rlabel metal1 215 -324 216 -323 1 q1
rlabel metal1 238 -324 239 -323 1 q2
rlabel m2contact 337 -382 337 -382 1 vdd
rlabel metal1 312 -372 313 -371 3 bl
rlabel metal1 361 -372 362 -371 7 blb
rlabel metal2 309 -364 309 -364 3 wl
rlabel metal1 325 -369 326 -368 5 q1
rlabel metal1 348 -369 349 -368 5 q2
rlabel m2contact 337 -346 337 -346 1 gnd
rlabel metal1 312 -321 313 -320 3 bl
rlabel metal1 361 -321 362 -320 7 blb
rlabel metal2 309 -328 309 -328 3 wl
rlabel metal1 325 -324 326 -323 1 q1
rlabel metal1 348 -324 349 -323 1 q2
rlabel metal1 257 -321 258 -320 3 bl
rlabel metal1 306 -321 307 -320 7 blb
rlabel metal2 254 -328 254 -328 3 wl
rlabel metal1 270 -324 271 -323 1 q1
rlabel metal1 293 -324 294 -323 1 q2
rlabel m2contact 447 -382 447 -382 1 vdd
rlabel metal1 422 -372 423 -371 3 bl
rlabel metal1 471 -372 472 -371 7 blb
rlabel metal2 419 -364 419 -364 3 wl
rlabel metal1 435 -369 436 -368 5 q1
rlabel metal1 458 -369 459 -368 5 q2
rlabel m2contact 392 -382 392 -382 1 vdd
rlabel metal1 367 -372 368 -371 3 bl
rlabel metal1 416 -372 417 -371 7 blb
rlabel metal2 364 -364 364 -364 3 wl
rlabel metal1 380 -369 381 -368 5 q1
rlabel metal1 403 -369 404 -368 5 q2
rlabel m2contact 447 -346 447 -346 1 gnd
rlabel metal1 422 -321 423 -320 3 bl
rlabel metal1 471 -321 472 -320 7 blb
rlabel metal2 419 -328 419 -328 3 wl
rlabel metal1 435 -324 436 -323 1 q1
rlabel metal1 458 -324 459 -323 1 q2
rlabel m2contact 392 -346 392 -346 1 gnd
rlabel metal1 367 -321 368 -320 3 bl
rlabel metal1 416 -321 417 -320 7 blb
rlabel metal2 364 -328 364 -328 3 wl
rlabel metal1 380 -324 381 -323 1 q1
rlabel metal1 403 -324 404 -323 1 q2
rlabel m2contact 612 -382 612 -382 1 vdd
rlabel metal1 587 -372 588 -371 3 bl
rlabel metal1 636 -372 637 -371 7 blb
rlabel metal2 584 -364 584 -364 3 wl
rlabel metal1 600 -369 601 -368 5 q1
rlabel metal1 623 -369 624 -368 5 q2
rlabel m2contact 557 -382 557 -382 1 vdd
rlabel metal1 532 -372 533 -371 3 bl
rlabel metal1 581 -372 582 -371 7 blb
rlabel metal2 529 -364 529 -364 3 wl
rlabel metal1 545 -369 546 -368 5 q1
rlabel metal1 568 -369 569 -368 5 q2
rlabel m2contact 502 -382 502 -382 1 vdd
rlabel metal1 477 -372 478 -371 3 bl
rlabel metal1 526 -372 527 -371 7 blb
rlabel metal2 474 -364 474 -364 3 wl
rlabel metal1 490 -369 491 -368 5 q1
rlabel metal1 513 -369 514 -368 5 q2
rlabel m2contact 612 -346 612 -346 1 gnd
rlabel metal1 587 -321 588 -320 3 bl
rlabel metal1 636 -321 637 -320 7 blb
rlabel metal2 584 -328 584 -328 3 wl
rlabel metal1 600 -324 601 -323 1 q1
rlabel metal1 623 -324 624 -323 1 q2
rlabel m2contact 557 -346 557 -346 1 gnd
rlabel metal1 532 -321 533 -320 3 bl
rlabel metal1 581 -321 582 -320 7 blb
rlabel metal2 529 -328 529 -328 3 wl
rlabel metal1 545 -324 546 -323 1 q1
rlabel metal1 568 -324 569 -323 1 q2
rlabel m2contact 502 -346 502 -346 1 gnd
rlabel metal1 477 -321 478 -320 3 bl
rlabel metal1 526 -321 527 -320 7 blb
rlabel metal2 474 -328 474 -328 3 wl
rlabel metal1 490 -324 491 -323 1 q1
rlabel metal1 513 -324 514 -323 1 q2
rlabel m2contact 282 -382 282 -382 1 vdd
rlabel m2contact 282 -346 282 -346 5 gnd
rlabel metal1 257 -372 258 -371 3 bl
rlabel metal1 306 -372 307 -371 7 blb
rlabel metal2 254 -364 254 -364 3 wl
rlabel metal1 270 -369 271 -368 5 q1
rlabel metal1 293 -369 294 -368 5 q2
rlabel m2contact 227 -310 227 -310 1 vdd
rlabel metal1 202 -300 203 -299 3 bl
rlabel metal1 251 -300 252 -299 7 blb
rlabel metal2 199 -292 199 -292 3 wl
rlabel metal1 215 -297 216 -296 5 q1
rlabel metal1 238 -297 239 -296 5 q2
rlabel m2contact 337 -310 337 -310 1 vdd
rlabel metal1 312 -300 313 -299 3 bl
rlabel metal1 361 -300 362 -299 7 blb
rlabel metal2 309 -292 309 -292 3 wl
rlabel metal1 325 -297 326 -296 5 q1
rlabel metal1 348 -297 349 -296 5 q2
rlabel m2contact 282 -310 282 -310 1 vdd
rlabel metal1 257 -300 258 -299 3 bl
rlabel metal1 306 -300 307 -299 7 blb
rlabel metal2 254 -292 254 -292 3 wl
rlabel metal1 270 -297 271 -296 5 q1
rlabel metal1 293 -297 294 -296 5 q2
rlabel m2contact 447 -310 447 -310 1 vdd
rlabel metal1 422 -300 423 -299 3 bl
rlabel metal1 471 -300 472 -299 7 blb
rlabel metal2 419 -292 419 -292 3 wl
rlabel metal1 435 -297 436 -296 5 q1
rlabel metal1 458 -297 459 -296 5 q2
rlabel m2contact 392 -310 392 -310 1 vdd
rlabel metal1 367 -300 368 -299 3 bl
rlabel metal1 416 -300 417 -299 7 blb
rlabel metal2 364 -292 364 -292 3 wl
rlabel metal1 380 -297 381 -296 5 q1
rlabel metal1 403 -297 404 -296 5 q2
rlabel m2contact 612 -310 612 -310 1 vdd
rlabel metal1 587 -300 588 -299 3 bl
rlabel metal1 636 -300 637 -299 7 blb
rlabel metal2 584 -292 584 -292 3 wl
rlabel metal1 600 -297 601 -296 5 q1
rlabel metal1 623 -297 624 -296 5 q2
rlabel m2contact 557 -310 557 -310 1 vdd
rlabel metal1 532 -300 533 -299 3 bl
rlabel metal1 581 -300 582 -299 7 blb
rlabel metal2 529 -292 529 -292 3 wl
rlabel metal1 545 -297 546 -296 5 q1
rlabel metal1 568 -297 569 -296 5 q2
rlabel m2contact 502 -310 502 -310 1 vdd
rlabel metal1 477 -300 478 -299 3 bl
rlabel metal1 526 -300 527 -299 7 blb
rlabel metal2 474 -292 474 -292 3 wl
rlabel metal1 490 -297 491 -296 5 q1
rlabel metal1 513 -297 514 -296 5 q2
rlabel m2contact 227 -274 227 -274 1 gnd
rlabel metal1 202 -249 203 -248 3 bl
rlabel metal1 251 -249 252 -248 7 blb
rlabel metal2 199 -256 199 -256 3 wl
rlabel metal1 215 -252 216 -251 1 q1
rlabel metal1 238 -252 239 -251 1 q2
rlabel m2contact 337 -274 337 -274 1 gnd
rlabel metal1 312 -249 313 -248 3 bl
rlabel metal1 361 -249 362 -248 7 blb
rlabel metal2 309 -256 309 -256 3 wl
rlabel metal1 325 -252 326 -251 1 q1
rlabel metal1 348 -252 349 -251 1 q2
rlabel metal1 257 -249 258 -248 3 bl
rlabel metal1 306 -249 307 -248 7 blb
rlabel metal2 254 -256 254 -256 3 wl
rlabel metal1 270 -252 271 -251 1 q1
rlabel metal1 293 -252 294 -251 1 q2
rlabel m2contact 447 -274 447 -274 1 gnd
rlabel metal1 422 -249 423 -248 3 bl
rlabel metal1 471 -249 472 -248 7 blb
rlabel metal2 419 -256 419 -256 3 wl
rlabel metal1 435 -252 436 -251 1 q1
rlabel metal1 458 -252 459 -251 1 q2
rlabel m2contact 392 -274 392 -274 1 gnd
rlabel metal1 367 -249 368 -248 3 bl
rlabel metal1 416 -249 417 -248 7 blb
rlabel metal2 364 -256 364 -256 3 wl
rlabel metal1 380 -252 381 -251 1 q1
rlabel metal1 403 -252 404 -251 1 q2
rlabel m2contact 612 -274 612 -274 1 gnd
rlabel metal1 587 -249 588 -248 3 bl
rlabel metal1 636 -249 637 -248 7 blb
rlabel metal2 584 -256 584 -256 3 wl
rlabel metal1 600 -252 601 -251 1 q1
rlabel metal1 623 -252 624 -251 1 q2
rlabel m2contact 557 -274 557 -274 1 gnd
rlabel metal1 532 -249 533 -248 3 bl
rlabel metal1 581 -249 582 -248 7 blb
rlabel metal2 529 -256 529 -256 3 wl
rlabel metal1 545 -252 546 -251 1 q1
rlabel metal1 568 -252 569 -251 1 q2
rlabel m2contact 502 -274 502 -274 1 gnd
rlabel metal1 477 -249 478 -248 3 bl
rlabel metal1 526 -249 527 -248 7 blb
rlabel metal2 474 -256 474 -256 3 wl
rlabel metal1 490 -252 491 -251 1 q1
rlabel metal1 513 -252 514 -251 1 q2
rlabel m2contact 282 -274 282 -274 5 gnd
rlabel m2contact 227 -238 227 -238 1 vdd
rlabel m2contact 337 -238 337 -238 1 vdd
rlabel m2contact 282 -238 282 -238 1 vdd
rlabel m2contact 447 -238 447 -238 1 vdd
rlabel m2contact 392 -238 392 -238 1 vdd
rlabel m2contact 612 -238 612 -238 1 vdd
rlabel m2contact 557 -238 557 -238 1 vdd
rlabel m2contact 502 -238 502 -238 1 vdd
<< end >>
