* SPICE3 file created from /home/swadesh/lab/magic/inverter/inverter.ext - technology: scmos
.lib /home/swadesh/cad/eda-technology/scn4m_subm/models/scn4m_cnrs_bsim3v1.lib nom

M1000 out in vdd vdd scmosp w=2u l=0.4u
+  ad=0p pd=0u as=0p ps=0u
M1001 out in gnd gnd scmosn w=1u l=0.4u
+  ad=0p pd=0u as=0p ps=0u
C0 vdd in 0.28fF
C1 in out 0.05fF
C2 vdd out 0.19fF
C3 out gnd 0.10fF
C4 in gnd 0.24fF
C5 vdd gnd 1.66fF

* TEST-BENCH *
.temp 27
.global vdd gnd


v0      vdd     gnd     dc      5
v1      in      gnd     pulse   0       5       1.5n    100p    100p    3n      6n
.tran 5p 15n
.control
run
plot v(out)+6 v(in)
.endc
.measure tran tdiff trig v(in) val=2.5 fall=1 targ v(out) val=2.5 rise=1
.measure tran tdiff trig v(in) val=2.5 rise=1 targ v(out) val=2.5 fall=1
.end
