magic
tech scmos
timestamp 1636288754
<< nwell >>
rect -13 -4 13 23
<< ntransistor >>
rect -1 -17 1 -13
<< ptransistor >>
rect -1 2 1 12
<< ndiffusion >>
rect -7 -17 -6 -13
rect -2 -17 -1 -13
rect 1 -17 2 -13
rect 6 -17 7 -13
<< pdiffusion >>
rect -7 11 -1 12
rect -7 3 -6 11
rect -2 3 -1 11
rect -7 2 -1 3
rect 1 11 7 12
rect 1 3 2 11
rect 6 3 7 11
rect 1 2 7 3
<< ndcontact >>
rect -6 -17 -2 -13
rect 2 -17 6 -13
<< pdcontact >>
rect -6 3 -2 11
rect 2 3 6 11
<< psubstratepcontact >>
rect -6 -25 -2 -21
rect 2 -25 6 -21
<< nsubstratencontact >>
rect -6 16 -2 20
rect 2 16 6 20
<< polysilicon >>
rect -1 12 1 14
rect -1 -5 1 2
rect -1 -13 1 -9
rect -1 -19 1 -17
<< polycontact >>
rect -3 -9 1 -5
<< metal1 >>
rect -7 16 -6 20
rect -2 16 2 20
rect 6 16 7 20
rect -6 11 -2 16
rect 6 3 7 11
rect 4 -13 7 3
rect 6 -17 7 -13
rect -6 -21 -2 -17
rect -7 -25 -6 -21
rect -2 -25 2 -21
rect 6 -25 7 -21
<< labels >>
rlabel metal1 0 18 0 18 5 vdd
rlabel metal1 0 -23 0 -23 1 gnd
rlabel metal1 5 -8 5 -8 1 out
rlabel polycontact -1 -7 -1 -7 1 in
<< end >>
