magic
tech scmos
timestamp 1635593005
<< nwell >>
rect 47 17 105 38
<< ntransistor >>
rect 56 5 60 8
rect 71 3 73 9
rect 79 3 81 9
rect 92 5 96 8
<< ptransistor >>
rect 67 24 73 27
rect 79 24 85 27
<< ndiffusion >>
rect 61 8 71 9
rect 55 5 56 8
rect 60 5 61 8
rect 68 4 71 8
rect 61 3 71 4
rect 73 8 79 9
rect 73 4 74 8
rect 78 4 79 8
rect 73 3 79 4
rect 81 8 91 9
rect 81 4 84 8
rect 91 5 92 8
rect 96 5 97 8
rect 81 3 91 4
<< pdiffusion >>
rect 66 24 67 27
rect 73 24 74 27
rect 78 24 79 27
rect 85 24 86 27
<< ndcontact >>
rect 51 4 55 8
rect 61 4 68 8
rect 74 4 78 8
rect 84 4 91 8
rect 97 4 101 8
<< pdcontact >>
rect 62 23 66 27
rect 74 24 78 28
rect 86 23 90 27
<< psubstratepcontact >>
rect 64 -5 68 -1
rect 84 -5 88 -1
<< nsubstratencontact >>
rect 62 31 66 35
rect 86 31 90 35
<< polysilicon >>
rect 67 27 73 29
rect 79 27 85 29
rect 67 22 73 24
rect 71 15 73 22
rect 56 8 60 13
rect 71 9 73 11
rect 79 22 85 24
rect 79 21 83 22
rect 79 9 81 17
rect 56 3 60 5
rect 92 8 96 13
rect 92 3 96 5
rect 71 1 73 3
rect 79 1 81 3
<< polycontact >>
rect 56 13 60 17
rect 69 11 73 15
rect 79 17 83 21
rect 92 13 96 17
<< metal1 >>
rect 50 8 53 38
rect 66 31 74 35
rect 78 31 86 35
rect 74 28 78 31
rect 63 21 66 23
rect 63 18 79 21
rect 63 8 66 18
rect 86 14 89 23
rect 73 11 89 14
rect 86 8 89 11
rect 99 8 102 38
rect 50 4 51 8
rect 101 4 102 8
rect 50 -8 53 4
rect 74 -1 78 4
rect 68 -5 74 -1
rect 78 -5 84 -1
rect 99 -8 102 4
<< m2contact >>
rect 74 31 78 35
rect 56 13 60 17
rect 92 13 96 17
rect 74 -5 78 -1
<< metal2 >>
rect 47 31 74 35
rect 78 31 105 35
rect 47 13 56 17
rect 60 13 92 17
rect 96 13 105 17
rect 47 -5 74 -1
rect 78 -5 105 -1
<< labels >>
rlabel m2contact 76 33 76 33 5 vdd
rlabel m2contact 76 -3 76 -3 1 gnd
rlabel metal1 51 22 52 23 3 bl
rlabel metal1 100 22 101 23 7 blb
rlabel metal2 48 15 48 15 3 wl
rlabel metal1 64 19 65 20 1 q1
rlabel metal1 87 19 88 20 1 q2
<< end >>
