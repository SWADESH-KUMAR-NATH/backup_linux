magic
tech scmos
timestamp 1627364388
<< nwell >>
rect 35 20 95 47
<< ntransistor >>
rect 47 9 49 14
rect 64 9 66 14
rect 81 9 83 14
<< ptransistor >>
rect 47 26 49 36
rect 64 26 66 36
rect 81 26 83 36
<< ndiffusion >>
rect 41 9 42 14
rect 46 9 47 14
rect 49 9 50 14
rect 54 9 55 14
rect 58 9 59 14
rect 63 9 64 14
rect 66 9 67 14
rect 71 9 72 14
rect 75 9 76 14
rect 80 9 81 14
rect 83 9 84 14
rect 88 9 89 14
<< pdiffusion >>
rect 41 35 47 36
rect 41 27 42 35
rect 46 27 47 35
rect 41 26 47 27
rect 49 35 55 36
rect 49 27 50 35
rect 54 27 55 35
rect 49 26 55 27
rect 58 35 64 36
rect 58 27 59 35
rect 63 27 64 35
rect 58 26 64 27
rect 66 35 72 36
rect 66 27 67 35
rect 71 27 72 35
rect 66 26 72 27
rect 75 35 81 36
rect 75 27 76 35
rect 80 27 81 35
rect 75 26 81 27
rect 83 35 89 36
rect 83 27 84 35
rect 88 27 89 35
rect 83 26 89 27
<< ndcontact >>
rect 42 9 46 14
rect 50 9 54 14
rect 59 9 63 14
rect 67 9 71 14
rect 76 9 80 14
rect 84 9 88 14
<< pdcontact >>
rect 42 27 46 35
rect 50 27 54 35
rect 59 27 63 35
rect 67 27 71 35
rect 76 27 80 35
rect 84 27 88 35
<< psubstratepcontact >>
rect 42 1 46 5
rect 50 1 54 5
rect 59 1 63 5
rect 67 1 71 5
rect 76 1 80 5
rect 84 1 88 5
<< nsubstratencontact >>
rect 42 40 46 44
rect 50 40 54 44
rect 59 40 63 44
rect 67 40 71 44
rect 76 40 80 44
rect 84 40 88 44
<< polysilicon >>
rect 47 36 49 38
rect 64 36 66 38
rect 81 36 83 38
rect 47 14 49 26
rect 64 14 66 26
rect 81 14 83 26
rect 47 7 49 9
rect 64 7 66 9
rect 81 7 83 9
<< polycontact >>
rect 43 18 47 22
rect 60 18 64 22
rect 77 18 81 22
<< metal1 >>
rect 39 44 90 45
rect 39 40 42 44
rect 46 40 50 44
rect 54 40 59 44
rect 63 40 67 44
rect 71 40 76 44
rect 80 40 84 44
rect 88 40 90 44
rect 39 39 90 40
rect 42 35 46 39
rect 59 35 63 39
rect 76 35 80 39
rect 50 22 54 27
rect 67 22 71 27
rect 84 22 88 27
rect 50 18 60 22
rect 67 18 77 22
rect 50 14 54 18
rect 67 14 71 18
rect 84 14 88 18
rect 42 6 46 9
rect 59 6 63 9
rect 76 6 80 9
rect 39 5 90 6
rect 39 1 42 5
rect 46 1 50 5
rect 54 1 59 5
rect 63 1 67 5
rect 71 1 76 5
rect 80 1 84 5
rect 88 1 90 5
rect 39 0 90 1
<< m2contact >>
rect 39 18 43 22
rect 84 18 88 22
<< metal2 >>
rect 43 18 84 22
<< labels >>
rlabel metal1 65 42 65 42 5 vdd
rlabel metal1 65 3 65 3 1 gnd
rlabel m2contact 86 20 86 20 1 out
<< end >>
