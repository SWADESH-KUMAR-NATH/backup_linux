magic
tech scmos
timestamp 1636469681
<< nwell >>
rect 0 -30 48 11
<< ntransistor >>
rect 11 -47 13 -38
rect 19 -47 21 -38
rect 35 -47 37 -38
<< ptransistor >>
rect 11 -24 13 0
rect 19 -24 21 -6
rect 27 -24 29 -6
rect 35 -24 37 0
<< ndiffusion >>
rect 6 -39 11 -38
rect 10 -46 11 -39
rect 6 -47 11 -46
rect 13 -39 19 -38
rect 13 -46 14 -39
rect 18 -46 19 -39
rect 13 -47 19 -46
rect 21 -39 26 -38
rect 21 -46 22 -39
rect 21 -47 26 -46
rect 30 -39 35 -38
rect 34 -46 35 -39
rect 30 -47 35 -46
rect 37 -39 42 -38
rect 37 -46 38 -39
rect 37 -47 42 -46
<< pdiffusion >>
rect 6 -1 11 0
rect 10 -23 11 -1
rect 6 -24 11 -23
rect 13 -1 18 0
rect 13 -23 14 -1
rect 30 -1 35 0
rect 18 -23 19 -6
rect 13 -24 19 -23
rect 21 -7 27 -6
rect 21 -23 22 -7
rect 26 -23 27 -7
rect 21 -24 27 -23
rect 29 -23 30 -6
rect 34 -23 35 -1
rect 29 -24 35 -23
rect 37 -1 42 0
rect 37 -23 38 -1
rect 37 -24 42 -23
<< ndcontact >>
rect 6 -46 10 -39
rect 14 -46 18 -39
rect 22 -46 26 -39
rect 30 -46 34 -39
rect 38 -46 42 -39
<< pdcontact >>
rect 6 -23 10 -1
rect 14 -23 18 -1
rect 22 -23 26 -7
rect 30 -23 34 -1
rect 38 -23 42 -1
<< psubstratepcontact >>
rect 38 -55 42 -51
<< nsubstratencontact >>
rect 14 4 18 8
rect 30 4 34 8
<< polysilicon >>
rect 11 1 37 3
rect 11 0 13 1
rect 35 0 37 1
rect 19 -6 21 -4
rect 27 -6 29 -4
rect 11 -26 13 -24
rect 19 -29 21 -24
rect 27 -26 29 -24
rect 14 -31 21 -29
rect 28 -30 29 -26
rect 14 -32 16 -31
rect 11 -36 12 -32
rect 24 -34 26 -30
rect 19 -36 26 -34
rect 11 -38 13 -36
rect 19 -38 21 -36
rect 35 -38 37 -24
rect 11 -49 13 -47
rect 19 -49 21 -47
rect 35 -61 37 -47
<< polycontact >>
rect 24 -30 28 -26
rect 12 -36 16 -32
rect 34 -65 38 -61
<< metal1 >>
rect 0 4 14 8
rect 18 4 30 8
rect 34 4 48 8
rect 22 -7 26 4
rect 14 -26 17 -23
rect 6 -29 24 -26
rect 6 -39 9 -29
rect 31 -33 34 -23
rect 16 -36 34 -33
rect 23 -39 26 -36
rect 14 -49 18 -46
rect 30 -49 34 -46
rect 14 -52 34 -49
rect 38 -51 42 -46
rect 0 -58 48 -55
rect 0 -65 34 -61
rect 38 -65 48 -61
<< m2contact >>
rect 6 -5 10 -1
rect 38 -5 42 -1
<< metal2 >>
rect 6 -1 9 8
rect 39 -1 42 8
rect 6 -65 9 -5
rect 39 -65 42 -5
<< labels >>
rlabel metal2 41 -28 41 -28 7 blb
rlabel metal2 7 -28 7 -28 3 bl
rlabel metal1 24 -63 24 -63 1 r_en
rlabel metal1 23 -57 23 -57 1 gnd
rlabel metal1 16 -27 16 -27 1 sa
rlabel metal1 32 -34 32 -34 1 sab
rlabel metal1 24 6 24 6 5 vdd
<< end >>
