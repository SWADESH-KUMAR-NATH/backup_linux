magic
tech scmos
timestamp 1636351123
<< nwell >>
rect -17 -7 17 20
<< ntransistor >>
rect -5 -20 -3 -14
rect 3 -20 5 -14
<< ptransistor >>
rect -5 0 -3 9
rect 3 0 5 9
<< ndiffusion >>
rect -11 -15 -5 -14
rect -11 -19 -10 -15
rect -6 -19 -5 -15
rect -11 -20 -5 -19
rect -3 -15 3 -14
rect -3 -19 -2 -15
rect 2 -19 3 -15
rect -3 -20 3 -19
rect 5 -15 11 -14
rect 5 -19 6 -15
rect 10 -19 11 -15
rect 5 -20 11 -19
<< pdiffusion >>
rect -11 8 -5 9
rect -11 1 -10 8
rect -6 1 -5 8
rect -11 0 -5 1
rect -3 8 3 9
rect -3 1 -2 8
rect 2 1 3 8
rect -3 0 3 1
rect 5 8 11 9
rect 5 1 6 8
rect 10 1 11 8
rect 5 0 11 1
<< ndcontact >>
rect -10 -19 -6 -15
rect -2 -19 2 -15
rect 6 -19 10 -15
<< pdcontact >>
rect -10 1 -6 8
rect -2 1 2 8
rect 6 1 10 8
<< psubstratepcontact >>
rect -2 -28 2 -24
<< nsubstratencontact >>
rect -2 13 2 17
<< polysilicon >>
rect -5 9 -3 11
rect 3 9 5 11
rect -5 -8 -3 0
rect 3 -8 5 0
rect -4 -12 -3 -8
rect 4 -12 5 -8
rect -5 -14 -3 -12
rect 3 -14 5 -12
rect -5 -22 -3 -20
rect 3 -22 5 -20
<< polycontact >>
rect -8 -12 -4 -8
rect 0 -12 4 -8
<< metal1 >>
rect -11 13 -2 17
rect 2 13 11 17
rect -2 8 2 13
rect 10 1 11 8
rect -10 -2 -7 1
rect 8 -2 11 1
rect -10 -5 11 -2
rect 8 -15 11 -5
rect 10 -19 11 -15
rect -10 -24 -6 -19
rect -11 -28 -2 -24
rect 2 -28 11 -24
<< labels >>
rlabel metal1 -8 -26 -8 -26 1 gnd
rlabel metal1 10 -5 10 -5 1 y
rlabel metal1 -8 15 -8 15 5 vdd
rlabel polycontact -6 -10 -6 -10 1 a
rlabel polycontact 2 -10 2 -10 1 b
<< end >>
