magic
tech scmos
timestamp 1635738960
<< nwell >>
rect -282 19 -261 21
rect -257 19 -223 21
rect -282 -13 -223 19
rect -282 -22 -279 -13
rect -271 -16 -235 -13
rect -271 -20 -260 -16
rect -251 -17 -235 -16
rect -246 -19 -235 -17
rect -245 -20 -235 -19
rect -271 -21 -263 -20
rect -261 -21 -253 -20
rect -244 -21 -235 -20
rect -271 -22 -250 -21
rect -242 -22 -235 -21
rect -227 -22 -223 -13
<< ntransistor >>
rect -271 43 -269 52
rect -263 43 -261 52
rect -245 43 -243 52
rect -237 43 -235 52
<< ndiffusion >>
rect -277 51 -271 52
rect -277 44 -276 51
rect -272 44 -271 51
rect -277 43 -271 44
rect -269 51 -263 52
rect -269 44 -268 51
rect -264 44 -263 51
rect -269 43 -263 44
rect -261 51 -255 52
rect -261 44 -260 51
rect -256 44 -255 51
rect -261 43 -255 44
rect -251 51 -245 52
rect -251 44 -250 51
rect -246 44 -245 51
rect -251 43 -245 44
rect -243 51 -237 52
rect -243 44 -242 51
rect -238 44 -237 51
rect -243 43 -237 44
rect -235 51 -229 52
rect -235 44 -234 51
rect -230 44 -229 51
rect -235 43 -229 44
<< ndcontact >>
rect -276 44 -272 51
rect -268 44 -264 51
rect -260 44 -256 51
rect -250 44 -246 51
rect -242 44 -238 51
rect -234 44 -230 51
<< psubstratepcontact >>
rect -276 35 -272 39
rect -268 35 -264 39
rect -259 35 -255 39
rect -251 35 -247 39
rect -242 35 -238 39
rect -234 35 -230 39
rect -268 -50 -264 -46
rect -242 -50 -238 -46
<< nsubstratencontact >>
rect -276 -3 -272 1
rect -268 -3 -264 1
rect -259 -3 -255 1
rect -251 -3 -247 1
rect -242 -3 -238 1
rect -234 -3 -230 1
<< polysilicon >>
rect -271 54 -268 56
rect -264 54 -261 56
rect -271 52 -269 54
rect -263 52 -261 54
rect -245 54 -242 56
rect -238 54 -235 56
rect -245 52 -243 54
rect -237 52 -235 54
rect -271 41 -269 43
rect -263 41 -261 43
rect -245 41 -243 43
rect -237 41 -235 43
<< polycontact >>
rect -268 54 -264 58
rect -242 54 -238 58
<< metal1 >>
rect -279 61 -256 64
rect -276 51 -273 61
rect -259 51 -256 61
rect -250 61 -227 64
rect -250 51 -247 61
rect -233 51 -230 61
rect -268 39 -264 44
rect -242 39 -238 44
rect -277 35 -276 39
rect -272 35 -268 39
rect -264 35 -259 39
rect -255 35 -251 39
rect -247 35 -242 39
rect -238 35 -234 39
rect -230 35 -229 39
rect -277 -3 -276 1
rect -272 -3 -268 1
rect -264 -3 -259 1
rect -255 -3 -251 1
rect -247 -3 -242 1
rect -238 -3 -234 1
rect -230 -3 -229 1
rect -270 -34 -240 -31
rect -277 -50 -268 -46
rect -264 -50 -242 -46
rect -238 -50 -229 -46
<< m2contact >>
rect -268 54 -264 58
rect -242 54 -238 58
rect -274 19 -270 23
rect -267 19 -263 23
rect -257 19 -253 23
rect -250 19 -246 23
rect -243 19 -239 23
rect -236 19 -232 23
rect -276 -25 -272 -21
rect -263 -28 -259 -24
rect -247 -28 -243 -24
rect -234 -25 -230 -21
rect -240 -34 -236 -30
<< metal2 >>
rect -267 23 -264 54
rect -242 23 -239 54
rect -275 19 -274 23
rect -232 19 -231 23
rect -275 -21 -272 19
rect -257 0 -254 19
rect -269 -3 -254 0
rect -269 -31 -266 -3
rect -249 -6 -246 19
rect -263 -9 -246 -6
rect -263 -24 -260 -9
rect -234 -21 -231 19
rect -255 -27 -247 -24
rect -255 -31 -252 -27
rect -283 -34 -252 -31
rect -249 -34 -240 -31
rect -249 -37 -246 -34
rect -283 -40 -246 -37
use nand  nand_2
timestamp 1633816195
transform -1 0 -266 0 1 -16
box -17 -34 17 20
use inv  inv_2
timestamp 1633895608
transform 1 0 -270 0 -1 17
box -13 -22 13 23
use nand  nand_3
timestamp 1633816195
transform 1 0 -240 0 1 -16
box -17 -34 17 20
use inv  inv_4
timestamp 1633895608
transform 1 0 -253 0 -1 17
box -13 -22 13 23
use inv  inv_3
timestamp 1633895608
transform -1 0 -236 0 -1 17
box -13 -22 13 23
<< labels >>
rlabel metal1 -253 -48 -253 -48 1 gnd
rlabel metal2 -281 -33 -281 -33 1 din
rlabel metal2 -281 -39 -281 -39 1 w_en
rlabel metal1 -277 62 -277 62 1 bl
rlabel metal1 -229 62 -229 62 1 blb
rlabel metal1 -253 36 -253 36 1 gnd
rlabel metal1 -253 -2 -253 -2 1 vdd
<< end >>
